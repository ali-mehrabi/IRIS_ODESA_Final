
module iris_auto_trainer
#(
parameter  p_sample_num = 75,
parameter  p_sample_len = 80,
parameter  p_spike_delay = 5,
parameter  p_pattern_delay = 5000,
parameter  p_epochs = 350
)
(
input         i_clk,
input         i_rst_n,
output        o_end_of_epochs,
output [4:1]  o_test_vector,
output [3:1]  o_label
);


parameter  p_test_len = (p_sample_num) * p_sample_len;


reg                                r_end_of_epochs;
reg   [2:0]                        r_state; 
reg   [$clog2(p_test_len-1):0]     r_address; 
reg   [7:1]                        r_data;
reg   [$clog2(p_pattern_delay):0]  r_counter;
reg   [$clog2(p_epochs):0]         r_epochs;
reg   [$clog2(p_spike_delay):0]    r_sp_counter;
wire  [7:1]                        r_ram[2249:0]; //[p_test_len-1:0];


assign o_test_vector = r_data[4:1];
assign o_label       = r_data[7:5];
assign o_end_of_epochs = r_end_of_epochs;

always @(posedge ~i_clk or negedge i_rst_n) 
begin 
if(!i_rst_n) 
  begin
    r_state   <= 0; 
	r_data    <= 0; 
	r_counter <= 0;
	r_address <= 0;
	r_epochs  <= 1;
	r_end_of_epochs <= 0;
	r_sp_counter <= 0;
  end
else 
   case(r_state) 
    0:begin 
	    if(r_counter < p_pattern_delay) 
		   r_counter <= r_counter+1;
		else 
		  begin
		    r_counter <= 0;
			r_state <= 1;
		  end
	  end
	1:begin
        r_data <= r_ram[r_address];
		r_state <= 2;
      end	
	2:begin
		r_data <= 0;
		if (r_sp_counter < p_spike_delay)
		   r_sp_counter <= r_sp_counter+1;
		else
		  begin
            r_sp_counter <= 0;
		    if(r_counter < p_sample_len - 1)
		      begin
		        r_counter <= r_counter+1;
			    r_address <= r_address+1;
				r_state <= 1;
		      end
		    else
		      begin
		        r_counter <= 0;
		  	    r_state <= 3;
		      end
		  end	  
	  end
	3:begin	
        //r_data <= 0;    
        if(r_counter < p_pattern_delay)
		  r_counter <= r_counter+1;
		else
		  begin
		    r_counter <= 0; 
		    if(r_address < (p_test_len-1)) 
              begin		
			    r_address <= r_address+1;
			    r_state <= 1;
			  end
			else
			  r_state <= 4;
		  end
	  end	  	
	4:begin
		if(r_epochs < p_epochs) 
		  begin
		    r_epochs <= r_epochs+1;
			r_address <= 0;
		    r_state <= 0;
		  end
		else
	      r_end_of_epochs <=1;
	  end		  
   endcase
end



// assign r_ram[0]= 7'h0;
// assign r_ram[1]= 7'h0;
// assign r_ram[2]= 7'h8;
// assign r_ram[3]= 7'h4;
// assign r_ram[4]= 7'h0;
// assign r_ram[5]= 7'h0;
// assign r_ram[6]= 7'h0;
// assign r_ram[7]= 7'h0;
// assign r_ram[8]= 7'h0;
// assign r_ram[9]= 7'h0;
// assign r_ram[10]= 7'h0;
// assign r_ram[11]= 7'h2;
// assign r_ram[12]= 7'h0;
// assign r_ram[13]= 7'h0;
// assign r_ram[14]= 7'h0;
// assign r_ram[15]= 7'h0;
// assign r_ram[16]= 7'h0;
// assign r_ram[17]= 7'h0;
// assign r_ram[18]= 7'h0;
// assign r_ram[19]= 7'h0;
// assign r_ram[20]= 7'h11;
// assign r_ram[21]= 7'h0;
// assign r_ram[22]= 7'h0;
// assign r_ram[23]= 7'h0;
// assign r_ram[24]= 7'h0;
// assign r_ram[25]= 7'h0;
// assign r_ram[26]= 7'h0;
// assign r_ram[27]= 7'h0;
// assign r_ram[28]= 7'h0;
// assign r_ram[29]= 7'h0;
// assign r_ram[30]= 7'h0;
// assign r_ram[31]= 7'h0;
// assign r_ram[32]= 7'h0;
// assign r_ram[33]= 7'h0;
// assign r_ram[34]= 7'h0;
// assign r_ram[35]= 7'h0;
// assign r_ram[36]= 7'h0;
// assign r_ram[37]= 7'h0;
// assign r_ram[38]= 7'h0;
// assign r_ram[39]= 7'h0;
// assign r_ram[40]= 7'h2;
// assign r_ram[41]= 7'h0;
// assign r_ram[42]= 7'h0;
// assign r_ram[43]= 7'h0;
// assign r_ram[44]= 7'h0;
// assign r_ram[45]= 7'h0;
// assign r_ram[46]= 7'h8;
// assign r_ram[47]= 7'h4;
// assign r_ram[48]= 7'h0;
// assign r_ram[49]= 7'h0;
// assign r_ram[50]= 7'h0;
// assign r_ram[51]= 7'h0;
// assign r_ram[52]= 7'h0;
// assign r_ram[53]= 7'h0;
// assign r_ram[54]= 7'h0;
// assign r_ram[55]= 7'h0;
// assign r_ram[56]= 7'h21;
// assign r_ram[57]= 7'h0;
// assign r_ram[58]= 7'h0;
// assign r_ram[59]= 7'h0;
// assign r_ram[60]= 7'h0;
// assign r_ram[61]= 7'h0;
// assign r_ram[62]= 7'h0;
// assign r_ram[63]= 7'h0;
// assign r_ram[64]= 7'h0;
// assign r_ram[65]= 7'h0;
// assign r_ram[66]= 7'h0;
// assign r_ram[67]= 7'h0;
// assign r_ram[68]= 7'h0;
// assign r_ram[69]= 7'h0;
// assign r_ram[70]= 7'h2;
// assign r_ram[71]= 7'h0;
// assign r_ram[72]= 7'h0;
// assign r_ram[73]= 7'h0;
// assign r_ram[74]= 7'h0;
// assign r_ram[75]= 7'h0;
// assign r_ram[76]= 7'h0;
// assign r_ram[77]= 7'h0;
// assign r_ram[78]= 7'h0;
// assign r_ram[79]= 7'h0;
// assign r_ram[80]= 7'h0;
// assign r_ram[81]= 7'h0;
// assign r_ram[82]= 7'h0;
// assign r_ram[83]= 7'h4;
// assign r_ram[84]= 7'h1;
// assign r_ram[85]= 7'h0;
// assign r_ram[86]= 7'h0;
// assign r_ram[87]= 7'h0;
// assign r_ram[88]= 7'h48;
// assign r_ram[89]= 7'h0;
// assign r_ram[90]= 7'h0;
// assign r_ram[91]= 7'h0;
// assign r_ram[92]= 7'h8;
// assign r_ram[93]= 7'h4;
// assign r_ram[94]= 7'h0;
// assign r_ram[95]= 7'h0;
// assign r_ram[96]= 7'h0;
// assign r_ram[97]= 7'h0;
// assign r_ram[98]= 7'h0;
// assign r_ram[99]= 7'h0;
// assign r_ram[100]= 7'h2;
// assign r_ram[101]= 7'h0;
// assign r_ram[102]= 7'h0;
// assign r_ram[103]= 7'h0;
// assign r_ram[104]= 7'h0;
// assign r_ram[105]= 7'h0;
// assign r_ram[106]= 7'h0;
// assign r_ram[107]= 7'h0;
// assign r_ram[108]= 7'h0;
// assign r_ram[109]= 7'h11;
// assign r_ram[110]= 7'h0;
// assign r_ram[111]= 7'h0;
// assign r_ram[112]= 7'h0;
// assign r_ram[113]= 7'h0;
// assign r_ram[114]= 7'h0;
// assign r_ram[115]= 7'h0;
// assign r_ram[116]= 7'h0;
// assign r_ram[117]= 7'h0;
// assign r_ram[118]= 7'h0;
// assign r_ram[119]= 7'h0;
// assign r_ram[120]= 7'h0;
// assign r_ram[121]= 7'h0;
// assign r_ram[122]= 7'h0;
// assign r_ram[123]= 7'h0;
// assign r_ram[124]= 7'h0;
// assign r_ram[125]= 7'h0;
// assign r_ram[126]= 7'h0;
// assign r_ram[127]= 7'h0;
// assign r_ram[128]= 7'h0;
// assign r_ram[129]= 7'h0;
// assign r_ram[130]= 7'h2;
// assign r_ram[131]= 7'h0;
// assign r_ram[132]= 7'h0;
// assign r_ram[133]= 7'h0;
// assign r_ram[134]= 7'h0;
// assign r_ram[135]= 7'h0;
// assign r_ram[136]= 7'h0;
// assign r_ram[137]= 7'hc;
// assign r_ram[138]= 7'h0;
// assign r_ram[139]= 7'h0;
// assign r_ram[140]= 7'h0;
// assign r_ram[141]= 7'h0;
// assign r_ram[142]= 7'h0;
// assign r_ram[143]= 7'h0;
// assign r_ram[144]= 7'h21;
// assign r_ram[145]= 7'h0;
// assign r_ram[146]= 7'h0;
// assign r_ram[147]= 7'h0;
// assign r_ram[148]= 7'h0;
// assign r_ram[149]= 7'h0;
// assign r_ram[150]= 7'h0;
// assign r_ram[151]= 7'h0;
// assign r_ram[152]= 7'h0;
// assign r_ram[153]= 7'h0;
// assign r_ram[154]= 7'h0;
// assign r_ram[155]= 7'h0;
// assign r_ram[156]= 7'h0;
// assign r_ram[157]= 7'h0;
// assign r_ram[158]= 7'h0;
// assign r_ram[159]= 7'h2;
// assign r_ram[160]= 7'h0;
// assign r_ram[161]= 7'h0;
// assign r_ram[162]= 7'h0;
// assign r_ram[163]= 7'h0;
// assign r_ram[164]= 7'h0;
// assign r_ram[165]= 7'h0;
// assign r_ram[166]= 7'h0;
// assign r_ram[167]= 7'h0;
// assign r_ram[168]= 7'h0;
// assign r_ram[169]= 7'h4;
// assign r_ram[170]= 7'h0;
// assign r_ram[171]= 7'h8;
// assign r_ram[172]= 7'h41;
// assign r_ram[173]= 7'h0;
// assign r_ram[174]= 7'h0;
// assign r_ram[175]= 7'h0;
// assign r_ram[176]= 7'h0;
// assign r_ram[177]= 7'h0;
// assign r_ram[178]= 7'h0;
// assign r_ram[179]= 7'h0;
// assign r_ram[180]= 7'h0;
// assign r_ram[181]= 7'h0;
// assign r_ram[182]= 7'h8;
// assign r_ram[183]= 7'h4;
// assign r_ram[184]= 7'h0;
// assign r_ram[185]= 7'h0;
// assign r_ram[186]= 7'h0;
// assign r_ram[187]= 7'h0;
// assign r_ram[188]= 7'h0;
// assign r_ram[189]= 7'h0;
// assign r_ram[190]= 7'h2;
// assign r_ram[191]= 7'h0;
// assign r_ram[192]= 7'h0;
// assign r_ram[193]= 7'h0;
// assign r_ram[194]= 7'h0;
// assign r_ram[195]= 7'h0;
// assign r_ram[196]= 7'h0;
// assign r_ram[197]= 7'h0;
// assign r_ram[198]= 7'h0;
// assign r_ram[199]= 7'h11;
// assign r_ram[200]= 7'h0;
// assign r_ram[201]= 7'h0;
// assign r_ram[202]= 7'h0;
// assign r_ram[203]= 7'h0;
// assign r_ram[204]= 7'h0;
// assign r_ram[205]= 7'h0;
// assign r_ram[206]= 7'h0;
// assign r_ram[207]= 7'h0;
// assign r_ram[208]= 7'h0;
// assign r_ram[209]= 7'h0;
// assign r_ram[210]= 7'h0;
// assign r_ram[211]= 7'h0;
// assign r_ram[212]= 7'h0;
// assign r_ram[213]= 7'h0;
// assign r_ram[214]= 7'h0;
// assign r_ram[215]= 7'h0;
// assign r_ram[216]= 7'h0;
// assign r_ram[217]= 7'h0;
// assign r_ram[218]= 7'h0;
// assign r_ram[219]= 7'h0;
// assign r_ram[220]= 7'h2;
// assign r_ram[221]= 7'h0;
// assign r_ram[222]= 7'h0;
// assign r_ram[223]= 7'h0;
// assign r_ram[224]= 7'h0;
// assign r_ram[225]= 7'h0;
// assign r_ram[226]= 7'h0;
// assign r_ram[227]= 7'h8;
// assign r_ram[228]= 7'h4;
// assign r_ram[229]= 7'h0;
// assign r_ram[230]= 7'h0;
// assign r_ram[231]= 7'h0;
// assign r_ram[232]= 7'h0;
// assign r_ram[233]= 7'h0;
// assign r_ram[234]= 7'h0;
// assign r_ram[235]= 7'h0;
// assign r_ram[236]= 7'h21;
// assign r_ram[237]= 7'h0;
// assign r_ram[238]= 7'h0;
// assign r_ram[239]= 7'h0;
// assign r_ram[240]= 7'h0;
// assign r_ram[241]= 7'h0;
// assign r_ram[242]= 7'h0;
// assign r_ram[243]= 7'h0;
// assign r_ram[244]= 7'h0;
// assign r_ram[245]= 7'h0;
// assign r_ram[246]= 7'h0;
// assign r_ram[247]= 7'h0;
// assign r_ram[248]= 7'h0;
// assign r_ram[249]= 7'h0;
// assign r_ram[250]= 7'h2;
// assign r_ram[251]= 7'h0;
// assign r_ram[252]= 7'h0;
// assign r_ram[253]= 7'h0;
// assign r_ram[254]= 7'h0;
// assign r_ram[255]= 7'h0;
// assign r_ram[256]= 7'h0;
// assign r_ram[257]= 7'h0;
// assign r_ram[258]= 7'h0;
// assign r_ram[259]= 7'h0;
// assign r_ram[260]= 7'h0;
// assign r_ram[261]= 7'h0;
// assign r_ram[262]= 7'h0;
// assign r_ram[263]= 7'hc;
// assign r_ram[264]= 7'h0;
// assign r_ram[265]= 7'h0;
// assign r_ram[266]= 7'h41;
// assign r_ram[267]= 7'h0;
// assign r_ram[268]= 7'h0;
// assign r_ram[269]= 7'h0;
// assign r_ram[270]= 7'h0;
// assign r_ram[271]= 7'h0;
// assign r_ram[272]= 7'h8;
// assign r_ram[273]= 7'h4;
// assign r_ram[274]= 7'h0;
// assign r_ram[275]= 7'h0;
// assign r_ram[276]= 7'h0;
// assign r_ram[277]= 7'h0;
// assign r_ram[278]= 7'h0;
// assign r_ram[279]= 7'h0;
// assign r_ram[280]= 7'h2;
// assign r_ram[281]= 7'h0;
// assign r_ram[282]= 7'h0;
// assign r_ram[283]= 7'h0;
// assign r_ram[284]= 7'h0;
// assign r_ram[285]= 7'h0;
// assign r_ram[286]= 7'h0;
// assign r_ram[287]= 7'h0;
// assign r_ram[288]= 7'h0;
// assign r_ram[289]= 7'h11;
// assign r_ram[290]= 7'h0;
// assign r_ram[291]= 7'h0;
// assign r_ram[292]= 7'h0;
// assign r_ram[293]= 7'h0;
// assign r_ram[294]= 7'h0;
// assign r_ram[295]= 7'h0;
// assign r_ram[296]= 7'h0;
// assign r_ram[297]= 7'h0;
// assign r_ram[298]= 7'h0;
// assign r_ram[299]= 7'h0;
// assign r_ram[300]= 7'h0;
// assign r_ram[301]= 7'h0;
// assign r_ram[302]= 7'h0;
// assign r_ram[303]= 7'h0;
// assign r_ram[304]= 7'h0;
// assign r_ram[305]= 7'h0;
// assign r_ram[306]= 7'h0;
// assign r_ram[307]= 7'h0;
// assign r_ram[308]= 7'h2;
// assign r_ram[309]= 7'h0;
// assign r_ram[310]= 7'h0;
// assign r_ram[311]= 7'h0;
// assign r_ram[312]= 7'h0;
// assign r_ram[313]= 7'h0;
// assign r_ram[314]= 7'h4;
// assign r_ram[315]= 7'h8;
// assign r_ram[316]= 7'h0;
// assign r_ram[317]= 7'h0;
// assign r_ram[318]= 7'h0;
// assign r_ram[319]= 7'h0;
// assign r_ram[320]= 7'h0;
// assign r_ram[321]= 7'h21;
// assign r_ram[322]= 7'h0;
// assign r_ram[323]= 7'h0;
// assign r_ram[324]= 7'h0;
// assign r_ram[325]= 7'h0;
// assign r_ram[326]= 7'h0;
// assign r_ram[327]= 7'h0;
// assign r_ram[328]= 7'h0;
// assign r_ram[329]= 7'h0;
// assign r_ram[330]= 7'h0;
// assign r_ram[331]= 7'h0;
// assign r_ram[332]= 7'h0;
// assign r_ram[333]= 7'h0;
// assign r_ram[334]= 7'h0;
// assign r_ram[335]= 7'h0;
// assign r_ram[336]= 7'h0;
// assign r_ram[337]= 7'h0;
// assign r_ram[338]= 7'h0;
// assign r_ram[339]= 7'h2;
// assign r_ram[340]= 7'h0;
// assign r_ram[341]= 7'h0;
// assign r_ram[342]= 7'h0;
// assign r_ram[343]= 7'h0;
// assign r_ram[344]= 7'h0;
// assign r_ram[345]= 7'h0;
// assign r_ram[346]= 7'h0;
// assign r_ram[347]= 7'h0;
// assign r_ram[348]= 7'h0;
// assign r_ram[349]= 7'h0;
// assign r_ram[350]= 7'h8;
// assign r_ram[351]= 7'h4;
// assign r_ram[352]= 7'h0;
// assign r_ram[353]= 7'h0;
// assign r_ram[354]= 7'h41;
// assign r_ram[355]= 7'h0;
// assign r_ram[356]= 7'h0;
// assign r_ram[357]= 7'h0;
// assign r_ram[358]= 7'h0;
// assign r_ram[359]= 7'h0;
// assign r_ram[360]= 7'h0;
// assign r_ram[361]= 7'h0;
// assign r_ram[362]= 7'h8;
// assign r_ram[363]= 7'h4;
// assign r_ram[364]= 7'h0;
// assign r_ram[365]= 7'h0;
// assign r_ram[366]= 7'h0;
// assign r_ram[367]= 7'h0;
// assign r_ram[368]= 7'h0;
// assign r_ram[369]= 7'h0;
// assign r_ram[370]= 7'h0;
// assign r_ram[371]= 7'h2;
// assign r_ram[372]= 7'h0;
// assign r_ram[373]= 7'h0;
// assign r_ram[374]= 7'h0;
// assign r_ram[375]= 7'h0;
// assign r_ram[376]= 7'h0;
// assign r_ram[377]= 7'h0;
// assign r_ram[378]= 7'h0;
// assign r_ram[379]= 7'h0;
// assign r_ram[380]= 7'h11;
// assign r_ram[381]= 7'h0;
// assign r_ram[382]= 7'h0;
// assign r_ram[383]= 7'h0;
// assign r_ram[384]= 7'h0;
// assign r_ram[385]= 7'h0;
// assign r_ram[386]= 7'h0;
// assign r_ram[387]= 7'h0;
// assign r_ram[388]= 7'h0;
// assign r_ram[389]= 7'h0;
// assign r_ram[390]= 7'h0;
// assign r_ram[391]= 7'h0;
// assign r_ram[392]= 7'h0;
// assign r_ram[393]= 7'h0;
// assign r_ram[394]= 7'h0;
// assign r_ram[395]= 7'h0;
// assign r_ram[396]= 7'h0;
// assign r_ram[397]= 7'h0;
// assign r_ram[398]= 7'h0;
// assign r_ram[399]= 7'h2;
// assign r_ram[400]= 7'h0;
// assign r_ram[401]= 7'h0;
// assign r_ram[402]= 7'h0;
// assign r_ram[403]= 7'h0;
// assign r_ram[404]= 7'h0;
// assign r_ram[405]= 7'h0;
// assign r_ram[406]= 7'h0;
// assign r_ram[407]= 7'hc;
// assign r_ram[408]= 7'h0;
// assign r_ram[409]= 7'h0;
// assign r_ram[410]= 7'h0;
// assign r_ram[411]= 7'h0;
// assign r_ram[412]= 7'h0;
// assign r_ram[413]= 7'h0;
// assign r_ram[414]= 7'h21;
// assign r_ram[415]= 7'h0;
// assign r_ram[416]= 7'h0;
// assign r_ram[417]= 7'h0;
// assign r_ram[418]= 7'h0;
// assign r_ram[419]= 7'h0;
// assign r_ram[420]= 7'h0;
// assign r_ram[421]= 7'h0;
// assign r_ram[422]= 7'h0;
// assign r_ram[423]= 7'h0;
// assign r_ram[424]= 7'h0;
// assign r_ram[425]= 7'h0;
// assign r_ram[426]= 7'h0;
// assign r_ram[427]= 7'h0;
// assign r_ram[428]= 7'h0;
// assign r_ram[429]= 7'h0;
// assign r_ram[430]= 7'h2;
// assign r_ram[431]= 7'h0;
// assign r_ram[432]= 7'h0;
// assign r_ram[433]= 7'h0;
// assign r_ram[434]= 7'h0;
// assign r_ram[435]= 7'h0;
// assign r_ram[436]= 7'h0;
// assign r_ram[437]= 7'h0;
// assign r_ram[438]= 7'h0;
// assign r_ram[439]= 7'h0;
// assign r_ram[440]= 7'h0;
// assign r_ram[441]= 7'h0;
// assign r_ram[442]= 7'h4;
// assign r_ram[443]= 7'h0;
// assign r_ram[444]= 7'h1;
// assign r_ram[445]= 7'h48;
// assign r_ram[446]= 7'h0;
// assign r_ram[447]= 7'h0;
// assign r_ram[448]= 7'h0;
// assign r_ram[449]= 7'h0;
// assign r_ram[450]= 7'h0;
// assign r_ram[451]= 7'h0;
// assign r_ram[452]= 7'h0;
// assign r_ram[453]= 7'h0;
// assign r_ram[454]= 7'hc;
// assign r_ram[455]= 7'h0;
// assign r_ram[456]= 7'h0;
// assign r_ram[457]= 7'h0;
// assign r_ram[458]= 7'h0;
// assign r_ram[459]= 7'h0;
// assign r_ram[460]= 7'h0;
// assign r_ram[461]= 7'h0;
// assign r_ram[462]= 7'h2;
// assign r_ram[463]= 7'h0;
// assign r_ram[464]= 7'h0;
// assign r_ram[465]= 7'h0;
// assign r_ram[466]= 7'h0;
// assign r_ram[467]= 7'h0;
// assign r_ram[468]= 7'h0;
// assign r_ram[469]= 7'h0;
// assign r_ram[470]= 7'h0;
// assign r_ram[471]= 7'h11;
// assign r_ram[472]= 7'h0;
// assign r_ram[473]= 7'h0;
// assign r_ram[474]= 7'h0;
// assign r_ram[475]= 7'h0;
// assign r_ram[476]= 7'h0;
// assign r_ram[477]= 7'h0;
// assign r_ram[478]= 7'h0;
// assign r_ram[479]= 7'h0;
// assign r_ram[480]= 7'h0;
// assign r_ram[481]= 7'h0;
// assign r_ram[482]= 7'h0;
// assign r_ram[483]= 7'h0;
// assign r_ram[484]= 7'h0;
// assign r_ram[485]= 7'h0;
// assign r_ram[486]= 7'h0;
// assign r_ram[487]= 7'h0;
// assign r_ram[488]= 7'h0;
// assign r_ram[489]= 7'h2;
// assign r_ram[490]= 7'h0;
// assign r_ram[491]= 7'h0;
// assign r_ram[492]= 7'h0;
// assign r_ram[493]= 7'h0;
// assign r_ram[494]= 7'h0;
// assign r_ram[495]= 7'h8;
// assign r_ram[496]= 7'h0;
// assign r_ram[497]= 7'h4;
// assign r_ram[498]= 7'h0;
// assign r_ram[499]= 7'h0;
// assign r_ram[500]= 7'h0;
// assign r_ram[501]= 7'h0;
// assign r_ram[502]= 7'h21;
// assign r_ram[503]= 7'h0;
// assign r_ram[504]= 7'h0;
// assign r_ram[505]= 7'h0;
// assign r_ram[506]= 7'h0;
// assign r_ram[507]= 7'h0;
// assign r_ram[508]= 7'h0;
// assign r_ram[509]= 7'h0;
// assign r_ram[510]= 7'h0;
// assign r_ram[511]= 7'h0;
// assign r_ram[512]= 7'h0;
// assign r_ram[513]= 7'h0;
// assign r_ram[514]= 7'h0;
// assign r_ram[515]= 7'h0;
// assign r_ram[516]= 7'h0;
// assign r_ram[517]= 7'h0;
// assign r_ram[518]= 7'h0;
// assign r_ram[519]= 7'h0;
// assign r_ram[520]= 7'h2;
// assign r_ram[521]= 7'h0;
// assign r_ram[522]= 7'h0;
// assign r_ram[523]= 7'h0;
// assign r_ram[524]= 7'h0;
// assign r_ram[525]= 7'h0;
// assign r_ram[526]= 7'h0;
// assign r_ram[527]= 7'h0;
// assign r_ram[528]= 7'h0;
// assign r_ram[529]= 7'h0;
// assign r_ram[530]= 7'h0;
// assign r_ram[531]= 7'h0;
// assign r_ram[532]= 7'h0;
// assign r_ram[533]= 7'h8;
// assign r_ram[534]= 7'h0;
// assign r_ram[535]= 7'h0;
// assign r_ram[536]= 7'h4;
// assign r_ram[537]= 7'h0;
// assign r_ram[538]= 7'h41;
// assign r_ram[539]= 7'h0;
// assign r_ram[540]= 7'h0;
// assign r_ram[541]= 7'h0;
// assign r_ram[542]= 7'h0;
// assign r_ram[543]= 7'hc;
// assign r_ram[544]= 7'h0;
// assign r_ram[545]= 7'h0;
// assign r_ram[546]= 7'h0;
// assign r_ram[547]= 7'h0;
// assign r_ram[548]= 7'h0;
// assign r_ram[549]= 7'h0;
// assign r_ram[550]= 7'h2;
// assign r_ram[551]= 7'h0;
// assign r_ram[552]= 7'h0;
// assign r_ram[553]= 7'h0;
// assign r_ram[554]= 7'h0;
// assign r_ram[555]= 7'h0;
// assign r_ram[556]= 7'h0;
// assign r_ram[557]= 7'h0;
// assign r_ram[558]= 7'h0;
// assign r_ram[559]= 7'h11;
// assign r_ram[560]= 7'h0;
// assign r_ram[561]= 7'h0;
// assign r_ram[562]= 7'h0;
// assign r_ram[563]= 7'h0;
// assign r_ram[564]= 7'h0;
// assign r_ram[565]= 7'h0;
// assign r_ram[566]= 7'h0;
// assign r_ram[567]= 7'h0;
// assign r_ram[568]= 7'h0;
// assign r_ram[569]= 7'h0;
// assign r_ram[570]= 7'h0;
// assign r_ram[571]= 7'h0;
// assign r_ram[572]= 7'h0;
// assign r_ram[573]= 7'h0;
// assign r_ram[574]= 7'h0;
// assign r_ram[575]= 7'h0;
// assign r_ram[576]= 7'h0;
// assign r_ram[577]= 7'h0;
// assign r_ram[578]= 7'h0;
// assign r_ram[579]= 7'h0;
// assign r_ram[580]= 7'h2;
// assign r_ram[581]= 7'h0;
// assign r_ram[582]= 7'h0;
// assign r_ram[583]= 7'h0;
// assign r_ram[584]= 7'h0;
// assign r_ram[585]= 7'h0;
// assign r_ram[586]= 7'h0;
// assign r_ram[587]= 7'h4;
// assign r_ram[588]= 7'h8;
// assign r_ram[589]= 7'h0;
// assign r_ram[590]= 7'h0;
// assign r_ram[591]= 7'h0;
// assign r_ram[592]= 7'h0;
// assign r_ram[593]= 7'h0;
// assign r_ram[594]= 7'h21;
// assign r_ram[595]= 7'h0;
// assign r_ram[596]= 7'h0;
// assign r_ram[597]= 7'h0;
// assign r_ram[598]= 7'h0;
// assign r_ram[599]= 7'h0;
// assign r_ram[600]= 7'h0;
// assign r_ram[601]= 7'h0;
// assign r_ram[602]= 7'h0;
// assign r_ram[603]= 7'h0;
// assign r_ram[604]= 7'h0;
// assign r_ram[605]= 7'h0;
// assign r_ram[606]= 7'h0;
// assign r_ram[607]= 7'h0;
// assign r_ram[608]= 7'h2;
// assign r_ram[609]= 7'h0;
// assign r_ram[610]= 7'h0;
// assign r_ram[611]= 7'h0;
// assign r_ram[612]= 7'h0;
// assign r_ram[613]= 7'h0;
// assign r_ram[614]= 7'h0;
// assign r_ram[615]= 7'h0;
// assign r_ram[616]= 7'h0;
// assign r_ram[617]= 7'h4;
// assign r_ram[618]= 7'h0;
// assign r_ram[619]= 7'h49;
// assign r_ram[620]= 7'h0;
// assign r_ram[621]= 7'h0;
// assign r_ram[622]= 7'h0;
// assign r_ram[623]= 7'h0;
// assign r_ram[624]= 7'h0;
// assign r_ram[625]= 7'h0;
// assign r_ram[626]= 7'h0;
// assign r_ram[627]= 7'h0;
// assign r_ram[628]= 7'h0;
// assign r_ram[629]= 7'h0;
// assign r_ram[630]= 7'h0;
// assign r_ram[631]= 7'h0;
// assign r_ram[632]= 7'h8;
// assign r_ram[633]= 7'h4;
// assign r_ram[634]= 7'h0;
// assign r_ram[635]= 7'h0;
// assign r_ram[636]= 7'h0;
// assign r_ram[637]= 7'h0;
// assign r_ram[638]= 7'h0;
// assign r_ram[639]= 7'h0;
// assign r_ram[640]= 7'h2;
// assign r_ram[641]= 7'h0;
// assign r_ram[642]= 7'h0;
// assign r_ram[643]= 7'h0;
// assign r_ram[644]= 7'h0;
// assign r_ram[645]= 7'h0;
// assign r_ram[646]= 7'h0;
// assign r_ram[647]= 7'h0;
// assign r_ram[648]= 7'h0;
// assign r_ram[649]= 7'h0;
// assign r_ram[650]= 7'h11;
// assign r_ram[651]= 7'h0;
// assign r_ram[652]= 7'h0;
// assign r_ram[653]= 7'h0;
// assign r_ram[654]= 7'h0;
// assign r_ram[655]= 7'h0;
// assign r_ram[656]= 7'h0;
// assign r_ram[657]= 7'h0;
// assign r_ram[658]= 7'h0;
// assign r_ram[659]= 7'h0;
// assign r_ram[660]= 7'h0;
// assign r_ram[661]= 7'h0;
// assign r_ram[662]= 7'h0;
// assign r_ram[663]= 7'h0;
// assign r_ram[664]= 7'h0;
// assign r_ram[665]= 7'h0;
// assign r_ram[666]= 7'h0;
// assign r_ram[667]= 7'h0;
// assign r_ram[668]= 7'h2;
// assign r_ram[669]= 7'h0;
// assign r_ram[670]= 7'h0;
// assign r_ram[671]= 7'hc;
// assign r_ram[672]= 7'h0;
// assign r_ram[673]= 7'h0;
// assign r_ram[674]= 7'h0;
// assign r_ram[675]= 7'h0;
// assign r_ram[676]= 7'h0;
// assign r_ram[677]= 7'h0;
// assign r_ram[678]= 7'h0;
// assign r_ram[679]= 7'h21;
// assign r_ram[680]= 7'h0;
// assign r_ram[681]= 7'h0;
// assign r_ram[682]= 7'h0;
// assign r_ram[683]= 7'h0;
// assign r_ram[684]= 7'h0;
// assign r_ram[685]= 7'h0;
// assign r_ram[686]= 7'h0;
// assign r_ram[687]= 7'h0;
// assign r_ram[688]= 7'h0;
// assign r_ram[689]= 7'h0;
// assign r_ram[690]= 7'h0;
// assign r_ram[691]= 7'h0;
// assign r_ram[692]= 7'h0;
// assign r_ram[693]= 7'h0;
// assign r_ram[694]= 7'h0;
// assign r_ram[695]= 7'h0;
// assign r_ram[696]= 7'h0;
// assign r_ram[697]= 7'h0;
// assign r_ram[698]= 7'h0;
// assign r_ram[699]= 7'h2;
// assign r_ram[700]= 7'h0;
// assign r_ram[701]= 7'h0;
// assign r_ram[702]= 7'h0;
// assign r_ram[703]= 7'h0;
// assign r_ram[704]= 7'h0;
// assign r_ram[705]= 7'h0;
// assign r_ram[706]= 7'h0;
// assign r_ram[707]= 7'h0;
// assign r_ram[708]= 7'h0;
// assign r_ram[709]= 7'h0;
// assign r_ram[710]= 7'h8;
// assign r_ram[711]= 7'h0;
// assign r_ram[712]= 7'h0;
// assign r_ram[713]= 7'h0;
// assign r_ram[714]= 7'h4;
// assign r_ram[715]= 7'h0;
// assign r_ram[716]= 7'h0;
// assign r_ram[717]= 7'h41;
// assign r_ram[718]= 7'h0;
// assign r_ram[719]= 7'h0;
// assign r_ram[720]= 7'h0;
// assign r_ram[721]= 7'h0;
// assign r_ram[722]= 7'h8;
// assign r_ram[723]= 7'h4;
// assign r_ram[724]= 7'h0;
// assign r_ram[725]= 7'h0;
// assign r_ram[726]= 7'h0;
// assign r_ram[727]= 7'h0;
// assign r_ram[728]= 7'h0;
// assign r_ram[729]= 7'h2;
// assign r_ram[730]= 7'h0;
// assign r_ram[731]= 7'h0;
// assign r_ram[732]= 7'h0;
// assign r_ram[733]= 7'h0;
// assign r_ram[734]= 7'h0;
// assign r_ram[735]= 7'h0;
// assign r_ram[736]= 7'h0;
// assign r_ram[737]= 7'h0;
// assign r_ram[738]= 7'h11;
// assign r_ram[739]= 7'h0;
// assign r_ram[740]= 7'h0;
// assign r_ram[741]= 7'h0;
// assign r_ram[742]= 7'h0;
// assign r_ram[743]= 7'h0;
// assign r_ram[744]= 7'h0;
// assign r_ram[745]= 7'h0;
// assign r_ram[746]= 7'h0;
// assign r_ram[747]= 7'h0;
// assign r_ram[748]= 7'h0;
// assign r_ram[749]= 7'h0;
// assign r_ram[750]= 7'h0;
// assign r_ram[751]= 7'h0;
// assign r_ram[752]= 7'h0;
// assign r_ram[753]= 7'h0;
// assign r_ram[754]= 7'h0;
// assign r_ram[755]= 7'h0;
// assign r_ram[756]= 7'h0;
// assign r_ram[757]= 7'h0;
// assign r_ram[758]= 7'h0;
// assign r_ram[759]= 7'h2;
// assign r_ram[760]= 7'h0;
// assign r_ram[761]= 7'h0;
// assign r_ram[762]= 7'h0;
// assign r_ram[763]= 7'h0;
// assign r_ram[764]= 7'h0;
// assign r_ram[765]= 7'h8;
// assign r_ram[766]= 7'h0;
// assign r_ram[767]= 7'h4;
// assign r_ram[768]= 7'h0;
// assign r_ram[769]= 7'h0;
// assign r_ram[770]= 7'h0;
// assign r_ram[771]= 7'h0;
// assign r_ram[772]= 7'h0;
// assign r_ram[773]= 7'h0;
// assign r_ram[774]= 7'h0;
// assign r_ram[775]= 7'h21;
// assign r_ram[776]= 7'h0;
// assign r_ram[777]= 7'h0;
// assign r_ram[778]= 7'h0;
// assign r_ram[779]= 7'h0;
// assign r_ram[780]= 7'h0;
// assign r_ram[781]= 7'h0;
// assign r_ram[782]= 7'h0;
// assign r_ram[783]= 7'h0;
// assign r_ram[784]= 7'h0;
// assign r_ram[785]= 7'h0;
// assign r_ram[786]= 7'h0;
// assign r_ram[787]= 7'h0;
// assign r_ram[788]= 7'h2;
// assign r_ram[789]= 7'h0;
// assign r_ram[790]= 7'h0;
// assign r_ram[791]= 7'h0;
// assign r_ram[792]= 7'h0;
// assign r_ram[793]= 7'h0;
// assign r_ram[794]= 7'h0;
// assign r_ram[795]= 7'h0;
// assign r_ram[796]= 7'h0;
// assign r_ram[797]= 7'h0;
// assign r_ram[798]= 7'h0;
// assign r_ram[799]= 7'h0;
// assign r_ram[800]= 7'h8;
// assign r_ram[801]= 7'h0;
// assign r_ram[802]= 7'h4;
// assign r_ram[803]= 7'h0;
// assign r_ram[804]= 7'h0;
// assign r_ram[805]= 7'h41;
// assign r_ram[806]= 7'h0;
// assign r_ram[807]= 7'h0;
// assign r_ram[808]= 7'h0;
// assign r_ram[809]= 7'h0;
// assign r_ram[810]= 7'h0;
// assign r_ram[811]= 7'h8;
// assign r_ram[812]= 7'h0;
// assign r_ram[813]= 7'h4;
// assign r_ram[814]= 7'h0;
// assign r_ram[815]= 7'h0;
// assign r_ram[816]= 7'h0;
// assign r_ram[817]= 7'h0;
// assign r_ram[818]= 7'h0;
// assign r_ram[819]= 7'h0;
// assign r_ram[820]= 7'h2;
// assign r_ram[821]= 7'h0;
// assign r_ram[822]= 7'h0;
// assign r_ram[823]= 7'h0;
// assign r_ram[824]= 7'h0;
// assign r_ram[825]= 7'h0;
// assign r_ram[826]= 7'h0;
// assign r_ram[827]= 7'h0;
// assign r_ram[828]= 7'h0;
// assign r_ram[829]= 7'h11;
// assign r_ram[830]= 7'h0;
// assign r_ram[831]= 7'h0;
// assign r_ram[832]= 7'h0;
// assign r_ram[833]= 7'h0;
// assign r_ram[834]= 7'h0;
// assign r_ram[835]= 7'h0;
// assign r_ram[836]= 7'h0;
// assign r_ram[837]= 7'h0;
// assign r_ram[838]= 7'h0;
// assign r_ram[839]= 7'h0;
// assign r_ram[840]= 7'h0;
// assign r_ram[841]= 7'h0;
// assign r_ram[842]= 7'h0;
// assign r_ram[843]= 7'h0;
// assign r_ram[844]= 7'h0;
// assign r_ram[845]= 7'h0;
// assign r_ram[846]= 7'h0;
// assign r_ram[847]= 7'h0;
// assign r_ram[848]= 7'h0;
// assign r_ram[849]= 7'h2;
// assign r_ram[850]= 7'h0;
// assign r_ram[851]= 7'h0;
// assign r_ram[852]= 7'h0;
// assign r_ram[853]= 7'h0;
// assign r_ram[854]= 7'h4;
// assign r_ram[855]= 7'h0;
// assign r_ram[856]= 7'h8;
// assign r_ram[857]= 7'h0;
// assign r_ram[858]= 7'h0;
// assign r_ram[859]= 7'h0;
// assign r_ram[860]= 7'h21;
// assign r_ram[861]= 7'h0;
// assign r_ram[862]= 7'h0;
// assign r_ram[863]= 7'h0;
// assign r_ram[864]= 7'h0;
// assign r_ram[865]= 7'h0;
// assign r_ram[866]= 7'h0;
// assign r_ram[867]= 7'h0;
// assign r_ram[868]= 7'h0;
// assign r_ram[869]= 7'h0;
// assign r_ram[870]= 7'h0;
// assign r_ram[871]= 7'h0;
// assign r_ram[872]= 7'h0;
// assign r_ram[873]= 7'h0;
// assign r_ram[874]= 7'h0;
// assign r_ram[875]= 7'h0;
// assign r_ram[876]= 7'h0;
// assign r_ram[877]= 7'h0;
// assign r_ram[878]= 7'h0;
// assign r_ram[879]= 7'h0;
// assign r_ram[880]= 7'h0;
// assign r_ram[881]= 7'h2;
// assign r_ram[882]= 7'h0;
// assign r_ram[883]= 7'h0;
// assign r_ram[884]= 7'h0;
// assign r_ram[885]= 7'h0;
// assign r_ram[886]= 7'h0;
// assign r_ram[887]= 7'h0;
// assign r_ram[888]= 7'h0;
// assign r_ram[889]= 7'h0;
// assign r_ram[890]= 7'h0;
// assign r_ram[891]= 7'h0;
// assign r_ram[892]= 7'h0;
// assign r_ram[893]= 7'h0;
// assign r_ram[894]= 7'h4;
// assign r_ram[895]= 7'h0;
// assign r_ram[896]= 7'h1;
// assign r_ram[897]= 7'h0;
// assign r_ram[898]= 7'h48;
// assign r_ram[899]= 7'h0;
// assign r_ram[900]= 7'h0;
// assign r_ram[901]= 7'h0;
// assign r_ram[902]= 7'h8;
// assign r_ram[903]= 7'h4;
// assign r_ram[904]= 7'h0;
// assign r_ram[905]= 7'h0;
// assign r_ram[906]= 7'h0;
// assign r_ram[907]= 7'h0;
// assign r_ram[908]= 7'h0;
// assign r_ram[909]= 7'h0;
// assign r_ram[910]= 7'h0;
// assign r_ram[911]= 7'h2;
// assign r_ram[912]= 7'h0;
// assign r_ram[913]= 7'h0;
// assign r_ram[914]= 7'h0;
// assign r_ram[915]= 7'h0;
// assign r_ram[916]= 7'h0;
// assign r_ram[917]= 7'h0;
// assign r_ram[918]= 7'h0;
// assign r_ram[919]= 7'h0;
// assign r_ram[920]= 7'h0;
// assign r_ram[921]= 7'h11;
// assign r_ram[922]= 7'h0;
// assign r_ram[923]= 7'h0;
// assign r_ram[924]= 7'h0;
// assign r_ram[925]= 7'h0;
// assign r_ram[926]= 7'h0;
// assign r_ram[927]= 7'h0;
// assign r_ram[928]= 7'h0;
// assign r_ram[929]= 7'h0;
// assign r_ram[930]= 7'h0;
// assign r_ram[931]= 7'h0;
// assign r_ram[932]= 7'h0;
// assign r_ram[933]= 7'h0;
// assign r_ram[934]= 7'h0;
// assign r_ram[935]= 7'h0;
// assign r_ram[936]= 7'h0;
// assign r_ram[937]= 7'h2;
// assign r_ram[938]= 7'h0;
// assign r_ram[939]= 7'h0;
// assign r_ram[940]= 7'h0;
// assign r_ram[941]= 7'h8;
// assign r_ram[942]= 7'h4;
// assign r_ram[943]= 7'h0;
// assign r_ram[944]= 7'h0;
// assign r_ram[945]= 7'h0;
// assign r_ram[946]= 7'h0;
// assign r_ram[947]= 7'h0;
// assign r_ram[948]= 7'h0;
// assign r_ram[949]= 7'h0;
// assign r_ram[950]= 7'h21;
// assign r_ram[951]= 7'h0;
// assign r_ram[952]= 7'h0;
// assign r_ram[953]= 7'h0;
// assign r_ram[954]= 7'h0;
// assign r_ram[955]= 7'h0;
// assign r_ram[956]= 7'h0;
// assign r_ram[957]= 7'h0;
// assign r_ram[958]= 7'h0;
// assign r_ram[959]= 7'h0;
// assign r_ram[960]= 7'h0;
// assign r_ram[961]= 7'h0;
// assign r_ram[962]= 7'h0;
// assign r_ram[963]= 7'h0;
// assign r_ram[964]= 7'h0;
// assign r_ram[965]= 7'h0;
// assign r_ram[966]= 7'h0;
// assign r_ram[967]= 7'h0;
// assign r_ram[968]= 7'h0;
// assign r_ram[969]= 7'h0;
// assign r_ram[970]= 7'h2;
// assign r_ram[971]= 7'h0;
// assign r_ram[972]= 7'h0;
// assign r_ram[973]= 7'h0;
// assign r_ram[974]= 7'h0;
// assign r_ram[975]= 7'h0;
// assign r_ram[976]= 7'h0;
// assign r_ram[977]= 7'h0;
// assign r_ram[978]= 7'h0;
// assign r_ram[979]= 7'h4;
// assign r_ram[980]= 7'h0;
// assign r_ram[981]= 7'h0;
// assign r_ram[982]= 7'h8;
// assign r_ram[983]= 7'h0;
// assign r_ram[984]= 7'h41;
// assign r_ram[985]= 7'h0;
// assign r_ram[986]= 7'h0;
// assign r_ram[987]= 7'h0;
// assign r_ram[988]= 7'h0;
// assign r_ram[989]= 7'h0;
// assign r_ram[990]= 7'h0;
// assign r_ram[991]= 7'h0;
// assign r_ram[992]= 7'h8;
// assign r_ram[993]= 7'h0;
// assign r_ram[994]= 7'h4;
// assign r_ram[995]= 7'h0;
// assign r_ram[996]= 7'h0;
// assign r_ram[997]= 7'h0;
// assign r_ram[998]= 7'h0;
// assign r_ram[999]= 7'h0;
// assign r_ram[1000]= 7'h2;
// assign r_ram[1001]= 7'h0;
// assign r_ram[1002]= 7'h0;
// assign r_ram[1003]= 7'h0;
// assign r_ram[1004]= 7'h0;
// assign r_ram[1005]= 7'h0;
// assign r_ram[1006]= 7'h0;
// assign r_ram[1007]= 7'h0;
// assign r_ram[1008]= 7'h0;
// assign r_ram[1009]= 7'h11;
// assign r_ram[1010]= 7'h0;
// assign r_ram[1011]= 7'h0;
// assign r_ram[1012]= 7'h0;
// assign r_ram[1013]= 7'h0;
// assign r_ram[1014]= 7'h0;
// assign r_ram[1015]= 7'h0;
// assign r_ram[1016]= 7'h0;
// assign r_ram[1017]= 7'h0;
// assign r_ram[1018]= 7'h0;
// assign r_ram[1019]= 7'h0;
// assign r_ram[1020]= 7'h0;
// assign r_ram[1021]= 7'h0;
// assign r_ram[1022]= 7'h0;
// assign r_ram[1023]= 7'h0;
// assign r_ram[1024]= 7'h0;
// assign r_ram[1025]= 7'h0;
// assign r_ram[1026]= 7'h0;
// assign r_ram[1027]= 7'h0;
// assign r_ram[1028]= 7'h0;
// assign r_ram[1029]= 7'h0;
// assign r_ram[1030]= 7'h2;
// assign r_ram[1031]= 7'h0;
// assign r_ram[1032]= 7'h0;
// assign r_ram[1033]= 7'h0;
// assign r_ram[1034]= 7'h0;
// assign r_ram[1035]= 7'h4;
// assign r_ram[1036]= 7'h0;
// assign r_ram[1037]= 7'h8;
// assign r_ram[1038]= 7'h0;
// assign r_ram[1039]= 7'h0;
// assign r_ram[1040]= 7'h0;
// assign r_ram[1041]= 7'h0;
// assign r_ram[1042]= 7'h21;
// assign r_ram[1043]= 7'h0;
// assign r_ram[1044]= 7'h0;
// assign r_ram[1045]= 7'h0;
// assign r_ram[1046]= 7'h0;
// assign r_ram[1047]= 7'h0;
// assign r_ram[1048]= 7'h0;
// assign r_ram[1049]= 7'h0;
// assign r_ram[1050]= 7'h0;
// assign r_ram[1051]= 7'h0;
// assign r_ram[1052]= 7'h0;
// assign r_ram[1053]= 7'h0;
// assign r_ram[1054]= 7'h0;
// assign r_ram[1055]= 7'h0;
// assign r_ram[1056]= 7'h0;
// assign r_ram[1057]= 7'h0;
// assign r_ram[1058]= 7'h0;
// assign r_ram[1059]= 7'h2;
// assign r_ram[1060]= 7'h0;
// assign r_ram[1061]= 7'h0;
// assign r_ram[1062]= 7'h0;
// assign r_ram[1063]= 7'h0;
// assign r_ram[1064]= 7'h0;
// assign r_ram[1065]= 7'h0;
// assign r_ram[1066]= 7'h0;
// assign r_ram[1067]= 7'h0;
// assign r_ram[1068]= 7'h0;
// assign r_ram[1069]= 7'h0;
// assign r_ram[1070]= 7'h4;
// assign r_ram[1071]= 7'h8;
// assign r_ram[1072]= 7'h0;
// assign r_ram[1073]= 7'h0;
// assign r_ram[1074]= 7'h41;
// assign r_ram[1075]= 7'h0;
// assign r_ram[1076]= 7'h0;
// assign r_ram[1077]= 7'h0;
// assign r_ram[1078]= 7'h0;
// assign r_ram[1079]= 7'h0;
// assign r_ram[1080]= 7'h0;
// assign r_ram[1081]= 7'h8;
// assign r_ram[1082]= 7'h0;
// assign r_ram[1083]= 7'h4;
// assign r_ram[1084]= 7'h0;
// assign r_ram[1085]= 7'h0;
// assign r_ram[1086]= 7'h0;
// assign r_ram[1087]= 7'h0;
// assign r_ram[1088]= 7'h0;
// assign r_ram[1089]= 7'h0;
// assign r_ram[1090]= 7'h2;
// assign r_ram[1091]= 7'h0;
// assign r_ram[1092]= 7'h0;
// assign r_ram[1093]= 7'h0;
// assign r_ram[1094]= 7'h0;
// assign r_ram[1095]= 7'h0;
// assign r_ram[1096]= 7'h0;
// assign r_ram[1097]= 7'h0;
// assign r_ram[1098]= 7'h0;
// assign r_ram[1099]= 7'h11;
// assign r_ram[1100]= 7'h0;
// assign r_ram[1101]= 7'h0;
// assign r_ram[1102]= 7'h0;
// assign r_ram[1103]= 7'h0;
// assign r_ram[1104]= 7'h0;
// assign r_ram[1105]= 7'h0;
// assign r_ram[1106]= 7'h0;
// assign r_ram[1107]= 7'h0;
// assign r_ram[1108]= 7'h0;
// assign r_ram[1109]= 7'h0;
// assign r_ram[1110]= 7'h0;
// assign r_ram[1111]= 7'h0;
// assign r_ram[1112]= 7'h0;
// assign r_ram[1113]= 7'h0;
// assign r_ram[1114]= 7'h0;
// assign r_ram[1115]= 7'h0;
// assign r_ram[1116]= 7'h0;
// assign r_ram[1117]= 7'h0;
// assign r_ram[1118]= 7'h2;
// assign r_ram[1119]= 7'h0;
// assign r_ram[1120]= 7'h0;
// assign r_ram[1121]= 7'h8;
// assign r_ram[1122]= 7'h0;
// assign r_ram[1123]= 7'h0;
// assign r_ram[1124]= 7'h4;
// assign r_ram[1125]= 7'h0;
// assign r_ram[1126]= 7'h0;
// assign r_ram[1127]= 7'h0;
// assign r_ram[1128]= 7'h0;
// assign r_ram[1129]= 7'h0;
// assign r_ram[1130]= 7'h0;
// assign r_ram[1131]= 7'h0;
// assign r_ram[1132]= 7'h0;
// assign r_ram[1133]= 7'h21;
// assign r_ram[1134]= 7'h0;
// assign r_ram[1135]= 7'h0;
// assign r_ram[1136]= 7'h0;
// assign r_ram[1137]= 7'h0;
// assign r_ram[1138]= 7'h0;
// assign r_ram[1139]= 7'h0;
// assign r_ram[1140]= 7'h0;
// assign r_ram[1141]= 7'h0;
// assign r_ram[1142]= 7'h0;
// assign r_ram[1143]= 7'h0;
// assign r_ram[1144]= 7'h0;
// assign r_ram[1145]= 7'h0;
// assign r_ram[1146]= 7'h0;
// assign r_ram[1147]= 7'h0;
// assign r_ram[1148]= 7'h0;
// assign r_ram[1149]= 7'h0;
// assign r_ram[1150]= 7'h2;
// assign r_ram[1151]= 7'h0;
// assign r_ram[1152]= 7'h0;
// assign r_ram[1153]= 7'h0;
// assign r_ram[1154]= 7'h0;
// assign r_ram[1155]= 7'h0;
// assign r_ram[1156]= 7'h0;
// assign r_ram[1157]= 7'h0;
// assign r_ram[1158]= 7'h0;
// assign r_ram[1159]= 7'h0;
// assign r_ram[1160]= 7'h0;
// assign r_ram[1161]= 7'h4;
// assign r_ram[1162]= 7'h0;
// assign r_ram[1163]= 7'h8;
// assign r_ram[1164]= 7'h0;
// assign r_ram[1165]= 7'h41;
// assign r_ram[1166]= 7'h0;
// assign r_ram[1167]= 7'h0;
// assign r_ram[1168]= 7'h0;
// assign r_ram[1169]= 7'h0;
// assign r_ram[1170]= 7'h0;
// assign r_ram[1171]= 7'h8;
// assign r_ram[1172]= 7'h4;
// assign r_ram[1173]= 7'h0;
// assign r_ram[1174]= 7'h0;
// assign r_ram[1175]= 7'h0;
// assign r_ram[1176]= 7'h0;
// assign r_ram[1177]= 7'h0;
// assign r_ram[1178]= 7'h0;
// assign r_ram[1179]= 7'h0;
// assign r_ram[1180]= 7'h2;
// assign r_ram[1181]= 7'h0;
// assign r_ram[1182]= 7'h0;
// assign r_ram[1183]= 7'h0;
// assign r_ram[1184]= 7'h0;
// assign r_ram[1185]= 7'h0;
// assign r_ram[1186]= 7'h0;
// assign r_ram[1187]= 7'h0;
// assign r_ram[1188]= 7'h11;
// assign r_ram[1189]= 7'h0;
// assign r_ram[1190]= 7'h0;
// assign r_ram[1191]= 7'h0;
// assign r_ram[1192]= 7'h0;
// assign r_ram[1193]= 7'h0;
// assign r_ram[1194]= 7'h0;
// assign r_ram[1195]= 7'h0;
// assign r_ram[1196]= 7'h0;
// assign r_ram[1197]= 7'h0;
// assign r_ram[1198]= 7'h0;
// assign r_ram[1199]= 7'h0;
// assign r_ram[1200]= 7'h0;
// assign r_ram[1201]= 7'h0;
// assign r_ram[1202]= 7'h0;
// assign r_ram[1203]= 7'h0;
// assign r_ram[1204]= 7'h0;
// assign r_ram[1205]= 7'h0;
// assign r_ram[1206]= 7'h0;
// assign r_ram[1207]= 7'h0;
// assign r_ram[1208]= 7'h0;
// assign r_ram[1209]= 7'h2;
// assign r_ram[1210]= 7'h0;
// assign r_ram[1211]= 7'h0;
// assign r_ram[1212]= 7'h0;
// assign r_ram[1213]= 7'h0;
// assign r_ram[1214]= 7'h0;
// assign r_ram[1215]= 7'h0;
// assign r_ram[1216]= 7'h8;
// assign r_ram[1217]= 7'h4;
// assign r_ram[1218]= 7'h0;
// assign r_ram[1219]= 7'h0;
// assign r_ram[1220]= 7'h0;
// assign r_ram[1221]= 7'h0;
// assign r_ram[1222]= 7'h0;
// assign r_ram[1223]= 7'h21;
// assign r_ram[1224]= 7'h0;
// assign r_ram[1225]= 7'h0;
// assign r_ram[1226]= 7'h0;
// assign r_ram[1227]= 7'h0;
// assign r_ram[1228]= 7'h0;
// assign r_ram[1229]= 7'h0;
// assign r_ram[1230]= 7'h0;
// assign r_ram[1231]= 7'h0;
// assign r_ram[1232]= 7'h0;
// assign r_ram[1233]= 7'h0;
// assign r_ram[1234]= 7'h0;
// assign r_ram[1235]= 7'h0;
// assign r_ram[1236]= 7'h0;
// assign r_ram[1237]= 7'h0;
// assign r_ram[1238]= 7'h2;
// assign r_ram[1239]= 7'h0;
// assign r_ram[1240]= 7'h0;
// assign r_ram[1241]= 7'h0;
// assign r_ram[1242]= 7'h0;
// assign r_ram[1243]= 7'h0;
// assign r_ram[1244]= 7'h0;
// assign r_ram[1245]= 7'h0;
// assign r_ram[1246]= 7'h0;
// assign r_ram[1247]= 7'h0;
// assign r_ram[1248]= 7'h0;
// assign r_ram[1249]= 7'h4;
// assign r_ram[1250]= 7'h0;
// assign r_ram[1251]= 7'h0;
// assign r_ram[1252]= 7'h49;
// assign r_ram[1253]= 7'h0;
// assign r_ram[1254]= 7'h0;
// assign r_ram[1255]= 7'h0;
// assign r_ram[1256]= 7'h0;
// assign r_ram[1257]= 7'h0;
// assign r_ram[1258]= 7'h0;
// assign r_ram[1259]= 7'h0;
// assign r_ram[1260]= 7'h0;
// assign r_ram[1261]= 7'h0;
// assign r_ram[1262]= 7'hc;
// assign r_ram[1263]= 7'h0;
// assign r_ram[1264]= 7'h0;
// assign r_ram[1265]= 7'h0;
// assign r_ram[1266]= 7'h0;
// assign r_ram[1267]= 7'h0;
// assign r_ram[1268]= 7'h0;
// assign r_ram[1269]= 7'h0;
// assign r_ram[1270]= 7'h0;
// assign r_ram[1271]= 7'h0;
// assign r_ram[1272]= 7'h2;
// assign r_ram[1273]= 7'h0;
// assign r_ram[1274]= 7'h0;
// assign r_ram[1275]= 7'h0;
// assign r_ram[1276]= 7'h0;
// assign r_ram[1277]= 7'h0;
// assign r_ram[1278]= 7'h0;
// assign r_ram[1279]= 7'h0;
// assign r_ram[1280]= 7'h0;
// assign r_ram[1281]= 7'h0;
// assign r_ram[1282]= 7'h11;
// assign r_ram[1283]= 7'h0;
// assign r_ram[1284]= 7'h0;
// assign r_ram[1285]= 7'h0;
// assign r_ram[1286]= 7'h0;
// assign r_ram[1287]= 7'h0;
// assign r_ram[1288]= 7'h0;
// assign r_ram[1289]= 7'h0;
// assign r_ram[1290]= 7'h0;
// assign r_ram[1291]= 7'h0;
// assign r_ram[1292]= 7'h0;
// assign r_ram[1293]= 7'h0;
// assign r_ram[1294]= 7'h0;
// assign r_ram[1295]= 7'h0;
// assign r_ram[1296]= 7'h0;
// assign r_ram[1297]= 7'h0;
// assign r_ram[1298]= 7'h0;
// assign r_ram[1299]= 7'h2;
// assign r_ram[1300]= 7'h0;
// assign r_ram[1301]= 7'h0;
// assign r_ram[1302]= 7'h0;
// assign r_ram[1303]= 7'h4;
// assign r_ram[1304]= 7'h0;
// assign r_ram[1305]= 7'h8;
// assign r_ram[1306]= 7'h0;
// assign r_ram[1307]= 7'h0;
// assign r_ram[1308]= 7'h0;
// assign r_ram[1309]= 7'h0;
// assign r_ram[1310]= 7'h0;
// assign r_ram[1311]= 7'h0;
// assign r_ram[1312]= 7'h21;
// assign r_ram[1313]= 7'h0;
// assign r_ram[1314]= 7'h0;
// assign r_ram[1315]= 7'h0;
// assign r_ram[1316]= 7'h0;
// assign r_ram[1317]= 7'h0;
// assign r_ram[1318]= 7'h0;
// assign r_ram[1319]= 7'h0;
// assign r_ram[1320]= 7'h0;
// assign r_ram[1321]= 7'h0;
// assign r_ram[1322]= 7'h0;
// assign r_ram[1323]= 7'h0;
// assign r_ram[1324]= 7'h0;
// assign r_ram[1325]= 7'h0;
// assign r_ram[1326]= 7'h0;
// assign r_ram[1327]= 7'h0;
// assign r_ram[1328]= 7'h0;
// assign r_ram[1329]= 7'h2;
// assign r_ram[1330]= 7'h0;
// assign r_ram[1331]= 7'h0;
// assign r_ram[1332]= 7'h0;
// assign r_ram[1333]= 7'h0;
// assign r_ram[1334]= 7'h0;
// assign r_ram[1335]= 7'h0;
// assign r_ram[1336]= 7'h0;
// assign r_ram[1337]= 7'h0;
// assign r_ram[1338]= 7'h0;
// assign r_ram[1339]= 7'h4;
// assign r_ram[1340]= 7'h0;
// assign r_ram[1341]= 7'h0;
// assign r_ram[1342]= 7'h1;
// assign r_ram[1343]= 7'h0;
// assign r_ram[1344]= 7'h0;
// assign r_ram[1345]= 7'h0;
// assign r_ram[1346]= 7'h0;
// assign r_ram[1347]= 7'h48;
// assign r_ram[1348]= 7'h0;
// assign r_ram[1349]= 7'h0;
// assign r_ram[1350]= 7'h0;
// assign r_ram[1351]= 7'h0;
// assign r_ram[1352]= 7'h0;
// assign r_ram[1353]= 7'h4;
// assign r_ram[1354]= 7'h8;
// assign r_ram[1355]= 7'h0;
// assign r_ram[1356]= 7'h0;
// assign r_ram[1357]= 7'h0;
// assign r_ram[1358]= 7'h0;
// assign r_ram[1359]= 7'h0;
// assign r_ram[1360]= 7'h0;
// assign r_ram[1361]= 7'h0;
// assign r_ram[1362]= 7'h0;
// assign r_ram[1363]= 7'h2;
// assign r_ram[1364]= 7'h0;
// assign r_ram[1365]= 7'h0;
// assign r_ram[1366]= 7'h0;
// assign r_ram[1367]= 7'h0;
// assign r_ram[1368]= 7'h0;
// assign r_ram[1369]= 7'h0;
// assign r_ram[1370]= 7'h0;
// assign r_ram[1371]= 7'h0;
// assign r_ram[1372]= 7'h11;
// assign r_ram[1373]= 7'h0;
// assign r_ram[1374]= 7'h0;
// assign r_ram[1375]= 7'h0;
// assign r_ram[1376]= 7'h0;
// assign r_ram[1377]= 7'h0;
// assign r_ram[1378]= 7'h0;
// assign r_ram[1379]= 7'h0;
// assign r_ram[1380]= 7'h0;
// assign r_ram[1381]= 7'h0;
// assign r_ram[1382]= 7'h0;
// assign r_ram[1383]= 7'h0;
// assign r_ram[1384]= 7'h0;
// assign r_ram[1385]= 7'h0;
// assign r_ram[1386]= 7'h0;
// assign r_ram[1387]= 7'h0;
// assign r_ram[1388]= 7'h0;
// assign r_ram[1389]= 7'h0;
// assign r_ram[1390]= 7'h2;
// assign r_ram[1391]= 7'h0;
// assign r_ram[1392]= 7'h0;
// assign r_ram[1393]= 7'h0;
// assign r_ram[1394]= 7'h0;
// assign r_ram[1395]= 7'h0;
// assign r_ram[1396]= 7'hc;
// assign r_ram[1397]= 7'h0;
// assign r_ram[1398]= 7'h0;
// assign r_ram[1399]= 7'h0;
// assign r_ram[1400]= 7'h0;
// assign r_ram[1401]= 7'h0;
// assign r_ram[1402]= 7'h0;
// assign r_ram[1403]= 7'h0;
// assign r_ram[1404]= 7'h0;
// assign r_ram[1405]= 7'h21;
// assign r_ram[1406]= 7'h0;
// assign r_ram[1407]= 7'h0;
// assign r_ram[1408]= 7'h0;
// assign r_ram[1409]= 7'h0;
// assign r_ram[1410]= 7'h0;
// assign r_ram[1411]= 7'h0;
// assign r_ram[1412]= 7'h0;
// assign r_ram[1413]= 7'h0;
// assign r_ram[1414]= 7'h0;
// assign r_ram[1415]= 7'h0;
// assign r_ram[1416]= 7'h0;
// assign r_ram[1417]= 7'h0;
// assign r_ram[1418]= 7'h0;
// assign r_ram[1419]= 7'h0;
// assign r_ram[1420]= 7'h2;
// assign r_ram[1421]= 7'h0;
// assign r_ram[1422]= 7'h0;
// assign r_ram[1423]= 7'h0;
// assign r_ram[1424]= 7'h0;
// assign r_ram[1425]= 7'h0;
// assign r_ram[1426]= 7'h0;
// assign r_ram[1427]= 7'h0;
// assign r_ram[1428]= 7'h0;
// assign r_ram[1429]= 7'h0;
// assign r_ram[1430]= 7'h4;
// assign r_ram[1431]= 7'h0;
// assign r_ram[1432]= 7'h0;
// assign r_ram[1433]= 7'h0;
// assign r_ram[1434]= 7'h1;
// assign r_ram[1435]= 7'h0;
// assign r_ram[1436]= 7'h48;
// assign r_ram[1437]= 7'h0;
// assign r_ram[1438]= 7'h0;
// assign r_ram[1439]= 7'h0;
// assign r_ram[1440]= 7'h0;
// assign r_ram[1441]= 7'h0;
// assign r_ram[1442]= 7'h0;
// assign r_ram[1443]= 7'h4;
// assign r_ram[1444]= 7'h8;
// assign r_ram[1445]= 7'h0;
// assign r_ram[1446]= 7'h0;
// assign r_ram[1447]= 7'h0;
// assign r_ram[1448]= 7'h0;
// assign r_ram[1449]= 7'h0;
// assign r_ram[1450]= 7'h0;
// assign r_ram[1451]= 7'h0;
// assign r_ram[1452]= 7'h2;
// assign r_ram[1453]= 7'h0;
// assign r_ram[1454]= 7'h0;
// assign r_ram[1455]= 7'h0;
// assign r_ram[1456]= 7'h0;
// assign r_ram[1457]= 7'h0;
// assign r_ram[1458]= 7'h0;
// assign r_ram[1459]= 7'h0;
// assign r_ram[1460]= 7'h0;
// assign r_ram[1461]= 7'h11;
// assign r_ram[1462]= 7'h0;
// assign r_ram[1463]= 7'h0;
// assign r_ram[1464]= 7'h0;
// assign r_ram[1465]= 7'h0;
// assign r_ram[1466]= 7'h0;
// assign r_ram[1467]= 7'h0;
// assign r_ram[1468]= 7'h0;
// assign r_ram[1469]= 7'h0;
// assign r_ram[1470]= 7'h0;
// assign r_ram[1471]= 7'h0;
// assign r_ram[1472]= 7'h0;
// assign r_ram[1473]= 7'h0;
// assign r_ram[1474]= 7'h0;
// assign r_ram[1475]= 7'h0;
// assign r_ram[1476]= 7'h0;
// assign r_ram[1477]= 7'h0;
// assign r_ram[1478]= 7'h0;
// assign r_ram[1479]= 7'h0;
// assign r_ram[1480]= 7'h2;
// assign r_ram[1481]= 7'h0;
// assign r_ram[1482]= 7'h0;
// assign r_ram[1483]= 7'h0;
// assign r_ram[1484]= 7'h0;
// assign r_ram[1485]= 7'h0;
// assign r_ram[1486]= 7'h0;
// assign r_ram[1487]= 7'hc;
// assign r_ram[1488]= 7'h0;
// assign r_ram[1489]= 7'h0;
// assign r_ram[1490]= 7'h0;
// assign r_ram[1491]= 7'h0;
// assign r_ram[1492]= 7'h21;
// assign r_ram[1493]= 7'h0;
// assign r_ram[1494]= 7'h0;
// assign r_ram[1495]= 7'h0;
// assign r_ram[1496]= 7'h0;
// assign r_ram[1497]= 7'h0;
// assign r_ram[1498]= 7'h0;
// assign r_ram[1499]= 7'h0;
// assign r_ram[1500]= 7'h0;
// assign r_ram[1501]= 7'h0;
// assign r_ram[1502]= 7'h0;
// assign r_ram[1503]= 7'h0;
// assign r_ram[1504]= 7'h0;
// assign r_ram[1505]= 7'h0;
// assign r_ram[1506]= 7'h0;
// assign r_ram[1507]= 7'h0;
// assign r_ram[1508]= 7'h0;
// assign r_ram[1509]= 7'h0;
// assign r_ram[1510]= 7'h2;
// assign r_ram[1511]= 7'h0;
// assign r_ram[1512]= 7'h0;
// assign r_ram[1513]= 7'h0;
// assign r_ram[1514]= 7'h0;
// assign r_ram[1515]= 7'h0;
// assign r_ram[1516]= 7'h0;
// assign r_ram[1517]= 7'h0;
// assign r_ram[1518]= 7'h0;
// assign r_ram[1519]= 7'h0;
// assign r_ram[1520]= 7'h8;
// assign r_ram[1521]= 7'h4;
// assign r_ram[1522]= 7'h0;
// assign r_ram[1523]= 7'h0;
// assign r_ram[1524]= 7'h41;
// assign r_ram[1525]= 7'h0;
// assign r_ram[1526]= 7'h0;
// assign r_ram[1527]= 7'h0;
// assign r_ram[1528]= 7'h0;
// assign r_ram[1529]= 7'h0;
// assign r_ram[1530]= 7'h0;
// assign r_ram[1531]= 7'h0;
// assign r_ram[1532]= 7'h0;
// assign r_ram[1533]= 7'hc;
// assign r_ram[1534]= 7'h0;
// assign r_ram[1535]= 7'h0;
// assign r_ram[1536]= 7'h0;
// assign r_ram[1537]= 7'h0;
// assign r_ram[1538]= 7'h0;
// assign r_ram[1539]= 7'h0;
// assign r_ram[1540]= 7'h0;
// assign r_ram[1541]= 7'h2;
// assign r_ram[1542]= 7'h0;
// assign r_ram[1543]= 7'h0;
// assign r_ram[1544]= 7'h0;
// assign r_ram[1545]= 7'h0;
// assign r_ram[1546]= 7'h0;
// assign r_ram[1547]= 7'h0;
// assign r_ram[1548]= 7'h0;
// assign r_ram[1549]= 7'h0;
// assign r_ram[1550]= 7'h11;
// assign r_ram[1551]= 7'h0;
// assign r_ram[1552]= 7'h0;
// assign r_ram[1553]= 7'h0;
// assign r_ram[1554]= 7'h0;
// assign r_ram[1555]= 7'h0;
// assign r_ram[1556]= 7'h0;
// assign r_ram[1557]= 7'h0;
// assign r_ram[1558]= 7'h0;
// assign r_ram[1559]= 7'h0;
// assign r_ram[1560]= 7'h0;
// assign r_ram[1561]= 7'h0;
// assign r_ram[1562]= 7'h0;
// assign r_ram[1563]= 7'h0;
// assign r_ram[1564]= 7'h0;
// assign r_ram[1565]= 7'h0;
// assign r_ram[1566]= 7'h0;
// assign r_ram[1567]= 7'h0;
// assign r_ram[1568]= 7'h0;
// assign r_ram[1569]= 7'h2;
// assign r_ram[1570]= 7'h0;
// assign r_ram[1571]= 7'h8;
// assign r_ram[1572]= 7'h0;
// assign r_ram[1573]= 7'h0;
// assign r_ram[1574]= 7'h0;
// assign r_ram[1575]= 7'h4;
// assign r_ram[1576]= 7'h0;
// assign r_ram[1577]= 7'h0;
// assign r_ram[1578]= 7'h0;
// assign r_ram[1579]= 7'h0;
// assign r_ram[1580]= 7'h0;
// assign r_ram[1581]= 7'h0;
// assign r_ram[1582]= 7'h21;
// assign r_ram[1583]= 7'h0;
// assign r_ram[1584]= 7'h0;
// assign r_ram[1585]= 7'h0;
// assign r_ram[1586]= 7'h0;
// assign r_ram[1587]= 7'h0;
// assign r_ram[1588]= 7'h0;
// assign r_ram[1589]= 7'h0;
// assign r_ram[1590]= 7'h0;
// assign r_ram[1591]= 7'h0;
// assign r_ram[1592]= 7'h0;
// assign r_ram[1593]= 7'h0;
// assign r_ram[1594]= 7'h0;
// assign r_ram[1595]= 7'h0;
// assign r_ram[1596]= 7'h0;
// assign r_ram[1597]= 7'h0;
// assign r_ram[1598]= 7'h0;
// assign r_ram[1599]= 7'h0;
// assign r_ram[1600]= 7'h0;
// assign r_ram[1601]= 7'h0;
// assign r_ram[1602]= 7'h2;
// assign r_ram[1603]= 7'h0;
// assign r_ram[1604]= 7'h0;
// assign r_ram[1605]= 7'h0;
// assign r_ram[1606]= 7'h0;
// assign r_ram[1607]= 7'h0;
// assign r_ram[1608]= 7'h0;
// assign r_ram[1609]= 7'h0;
// assign r_ram[1610]= 7'h0;
// assign r_ram[1611]= 7'h0;
// assign r_ram[1612]= 7'h0;
// assign r_ram[1613]= 7'h0;
// assign r_ram[1614]= 7'h0;
// assign r_ram[1615]= 7'h8;
// assign r_ram[1616]= 7'h4;
// assign r_ram[1617]= 7'h0;
// assign r_ram[1618]= 7'h41;
// assign r_ram[1619]= 7'h0;
// assign r_ram[1620]= 7'h0;
// assign r_ram[1621]= 7'h0;
// assign r_ram[1622]= 7'h0;
// assign r_ram[1623]= 7'h8;
// assign r_ram[1624]= 7'h4;
// assign r_ram[1625]= 7'h0;
// assign r_ram[1626]= 7'h0;
// assign r_ram[1627]= 7'h0;
// assign r_ram[1628]= 7'h0;
// assign r_ram[1629]= 7'h0;
// assign r_ram[1630]= 7'h0;
// assign r_ram[1631]= 7'h0;
// assign r_ram[1632]= 7'h2;
// assign r_ram[1633]= 7'h0;
// assign r_ram[1634]= 7'h0;
// assign r_ram[1635]= 7'h0;
// assign r_ram[1636]= 7'h0;
// assign r_ram[1637]= 7'h0;
// assign r_ram[1638]= 7'h0;
// assign r_ram[1639]= 7'h0;
// assign r_ram[1640]= 7'h0;
// assign r_ram[1641]= 7'h0;
// assign r_ram[1642]= 7'h11;
// assign r_ram[1643]= 7'h0;
// assign r_ram[1644]= 7'h0;
// assign r_ram[1645]= 7'h0;
// assign r_ram[1646]= 7'h0;
// assign r_ram[1647]= 7'h0;
// assign r_ram[1648]= 7'h0;
// assign r_ram[1649]= 7'h0;
// assign r_ram[1650]= 7'h0;
// assign r_ram[1651]= 7'h0;
// assign r_ram[1652]= 7'h0;
// assign r_ram[1653]= 7'h0;
// assign r_ram[1654]= 7'h0;
// assign r_ram[1655]= 7'h0;
// assign r_ram[1656]= 7'h0;
// assign r_ram[1657]= 7'h0;
// assign r_ram[1658]= 7'h2;
// assign r_ram[1659]= 7'h0;
// assign r_ram[1660]= 7'h0;
// assign r_ram[1661]= 7'h0;
// assign r_ram[1662]= 7'h0;
// assign r_ram[1663]= 7'h0;
// assign r_ram[1664]= 7'h0;
// assign r_ram[1665]= 7'h0;
// assign r_ram[1666]= 7'h0;
// assign r_ram[1667]= 7'hc;
// assign r_ram[1668]= 7'h0;
// assign r_ram[1669]= 7'h0;
// assign r_ram[1670]= 7'h0;
// assign r_ram[1671]= 7'h0;
// assign r_ram[1672]= 7'h0;
// assign r_ram[1673]= 7'h21;
// assign r_ram[1674]= 7'h0;
// assign r_ram[1675]= 7'h0;
// assign r_ram[1676]= 7'h0;
// assign r_ram[1677]= 7'h0;
// assign r_ram[1678]= 7'h0;
// assign r_ram[1679]= 7'h0;
// assign r_ram[1680]= 7'h0;
// assign r_ram[1681]= 7'h0;
// assign r_ram[1682]= 7'h0;
// assign r_ram[1683]= 7'h0;
// assign r_ram[1684]= 7'h0;
// assign r_ram[1685]= 7'h0;
// assign r_ram[1686]= 7'h0;
// assign r_ram[1687]= 7'h0;
// assign r_ram[1688]= 7'h2;
// assign r_ram[1689]= 7'h0;
// assign r_ram[1690]= 7'h0;
// assign r_ram[1691]= 7'h0;
// assign r_ram[1692]= 7'h0;
// assign r_ram[1693]= 7'h0;
// assign r_ram[1694]= 7'h0;
// assign r_ram[1695]= 7'h0;
// assign r_ram[1696]= 7'h0;
// assign r_ram[1697]= 7'h0;
// assign r_ram[1698]= 7'h0;
// assign r_ram[1699]= 7'h0;
// assign r_ram[1700]= 7'h0;
// assign r_ram[1701]= 7'h0;
// assign r_ram[1702]= 7'h0;
// assign r_ram[1703]= 7'h0;
// assign r_ram[1704]= 7'h0;
// assign r_ram[1705]= 7'h0;
// assign r_ram[1706]= 7'h8;
// assign r_ram[1707]= 7'h4;
// assign r_ram[1708]= 7'h41;
// assign r_ram[1709]= 7'h0;
// assign r_ram[1710]= 7'h0;
// assign r_ram[1711]= 7'h0;
// assign r_ram[1712]= 7'h0;
// assign r_ram[1713]= 7'hc;
// assign r_ram[1714]= 7'h0;
// assign r_ram[1715]= 7'h0;
// assign r_ram[1716]= 7'h0;
// assign r_ram[1717]= 7'h0;
// assign r_ram[1718]= 7'h0;
// assign r_ram[1719]= 7'h0;
// assign r_ram[1720]= 7'h0;
// assign r_ram[1721]= 7'h0;
// assign r_ram[1722]= 7'h2;
// assign r_ram[1723]= 7'h0;
// assign r_ram[1724]= 7'h0;
// assign r_ram[1725]= 7'h0;
// assign r_ram[1726]= 7'h0;
// assign r_ram[1727]= 7'h0;
// assign r_ram[1728]= 7'h0;
// assign r_ram[1729]= 7'h0;
// assign r_ram[1730]= 7'h11;
// assign r_ram[1731]= 7'h0;
// assign r_ram[1732]= 7'h0;
// assign r_ram[1733]= 7'h0;
// assign r_ram[1734]= 7'h0;
// assign r_ram[1735]= 7'h0;
// assign r_ram[1736]= 7'h0;
// assign r_ram[1737]= 7'h0;
// assign r_ram[1738]= 7'h0;
// assign r_ram[1739]= 7'h0;
// assign r_ram[1740]= 7'h0;
// assign r_ram[1741]= 7'h0;
// assign r_ram[1742]= 7'h0;
// assign r_ram[1743]= 7'h0;
// assign r_ram[1744]= 7'h0;
// assign r_ram[1745]= 7'h0;
// assign r_ram[1746]= 7'h0;
// assign r_ram[1747]= 7'h0;
// assign r_ram[1748]= 7'h2;
// assign r_ram[1749]= 7'h0;
// assign r_ram[1750]= 7'h0;
// assign r_ram[1751]= 7'h0;
// assign r_ram[1752]= 7'h8;
// assign r_ram[1753]= 7'h0;
// assign r_ram[1754]= 7'h4;
// assign r_ram[1755]= 7'h0;
// assign r_ram[1756]= 7'h0;
// assign r_ram[1757]= 7'h0;
// assign r_ram[1758]= 7'h0;
// assign r_ram[1759]= 7'h0;
// assign r_ram[1760]= 7'h0;
// assign r_ram[1761]= 7'h0;
// assign r_ram[1762]= 7'h21;
// assign r_ram[1763]= 7'h0;
// assign r_ram[1764]= 7'h0;
// assign r_ram[1765]= 7'h0;
// assign r_ram[1766]= 7'h0;
// assign r_ram[1767]= 7'h0;
// assign r_ram[1768]= 7'h0;
// assign r_ram[1769]= 7'h0;
// assign r_ram[1770]= 7'h0;
// assign r_ram[1771]= 7'h0;
// assign r_ram[1772]= 7'h0;
// assign r_ram[1773]= 7'h0;
// assign r_ram[1774]= 7'h0;
// assign r_ram[1775]= 7'h0;
// assign r_ram[1776]= 7'h0;
// assign r_ram[1777]= 7'h0;
// assign r_ram[1778]= 7'h2;
// assign r_ram[1779]= 7'h0;
// assign r_ram[1780]= 7'h0;
// assign r_ram[1781]= 7'h0;
// assign r_ram[1782]= 7'h0;
// assign r_ram[1783]= 7'h0;
// assign r_ram[1784]= 7'h0;
// assign r_ram[1785]= 7'h0;
// assign r_ram[1786]= 7'h0;
// assign r_ram[1787]= 7'h8;
// assign r_ram[1788]= 7'h0;
// assign r_ram[1789]= 7'h4;
// assign r_ram[1790]= 7'h0;
// assign r_ram[1791]= 7'h0;
// assign r_ram[1792]= 7'h0;
// assign r_ram[1793]= 7'h41;
// assign r_ram[1794]= 7'h0;
// assign r_ram[1795]= 7'h0;
// assign r_ram[1796]= 7'h0;
// assign r_ram[1797]= 7'h0;
// assign r_ram[1798]= 7'h0;
// assign r_ram[1799]= 7'h0;
// assign r_ram[1800]= 7'h0;
// assign r_ram[1801]= 7'h0;
// assign r_ram[1802]= 7'h8;
// assign r_ram[1803]= 7'h0;
// assign r_ram[1804]= 7'h4;
// assign r_ram[1805]= 7'h0;
// assign r_ram[1806]= 7'h0;
// assign r_ram[1807]= 7'h0;
// assign r_ram[1808]= 7'h0;
// assign r_ram[1809]= 7'h0;
// assign r_ram[1810]= 7'h2;
// assign r_ram[1811]= 7'h0;
// assign r_ram[1812]= 7'h0;
// assign r_ram[1813]= 7'h0;
// assign r_ram[1814]= 7'h0;
// assign r_ram[1815]= 7'h0;
// assign r_ram[1816]= 7'h0;
// assign r_ram[1817]= 7'h0;
// assign r_ram[1818]= 7'h0;
// assign r_ram[1819]= 7'h0;
// assign r_ram[1820]= 7'h0;
// assign r_ram[1821]= 7'h11;
// assign r_ram[1822]= 7'h0;
// assign r_ram[1823]= 7'h0;
// assign r_ram[1824]= 7'h0;
// assign r_ram[1825]= 7'h0;
// assign r_ram[1826]= 7'h0;
// assign r_ram[1827]= 7'h0;
// assign r_ram[1828]= 7'h0;
// assign r_ram[1829]= 7'h0;
// assign r_ram[1830]= 7'h0;
// assign r_ram[1831]= 7'h0;
// assign r_ram[1832]= 7'h0;
// assign r_ram[1833]= 7'h0;
// assign r_ram[1834]= 7'h0;
// assign r_ram[1835]= 7'h0;
// assign r_ram[1836]= 7'h0;
// assign r_ram[1837]= 7'h0;
// assign r_ram[1838]= 7'h0;
// assign r_ram[1839]= 7'h0;
// assign r_ram[1840]= 7'h2;
// assign r_ram[1841]= 7'h0;
// assign r_ram[1842]= 7'h0;
// assign r_ram[1843]= 7'h0;
// assign r_ram[1844]= 7'h0;
// assign r_ram[1845]= 7'h0;
// assign r_ram[1846]= 7'h0;
// assign r_ram[1847]= 7'h0;
// assign r_ram[1848]= 7'h4;
// assign r_ram[1849]= 7'h0;
// assign r_ram[1850]= 7'h8;
// assign r_ram[1851]= 7'h0;
// assign r_ram[1852]= 7'h21;
// assign r_ram[1853]= 7'h0;
// assign r_ram[1854]= 7'h0;
// assign r_ram[1855]= 7'h0;
// assign r_ram[1856]= 7'h0;
// assign r_ram[1857]= 7'h0;
// assign r_ram[1858]= 7'h0;
// assign r_ram[1859]= 7'h0;
// assign r_ram[1860]= 7'h0;
// assign r_ram[1861]= 7'h0;
// assign r_ram[1862]= 7'h0;
// assign r_ram[1863]= 7'h0;
// assign r_ram[1864]= 7'h0;
// assign r_ram[1865]= 7'h0;
// assign r_ram[1866]= 7'h0;
// assign r_ram[1867]= 7'h0;
// assign r_ram[1868]= 7'h0;
// assign r_ram[1869]= 7'h0;
// assign r_ram[1870]= 7'h2;
// assign r_ram[1871]= 7'h0;
// assign r_ram[1872]= 7'h0;
// assign r_ram[1873]= 7'h0;
// assign r_ram[1874]= 7'h0;
// assign r_ram[1875]= 7'h0;
// assign r_ram[1876]= 7'h0;
// assign r_ram[1877]= 7'h0;
// assign r_ram[1878]= 7'h0;
// assign r_ram[1879]= 7'h0;
// assign r_ram[1880]= 7'h0;
// assign r_ram[1881]= 7'h0;
// assign r_ram[1882]= 7'h4;
// assign r_ram[1883]= 7'h0;
// assign r_ram[1884]= 7'h0;
// assign r_ram[1885]= 7'h0;
// assign r_ram[1886]= 7'h49;
// assign r_ram[1887]= 7'h0;
// assign r_ram[1888]= 7'h0;
// assign r_ram[1889]= 7'h0;
// assign r_ram[1890]= 7'h0;
// assign r_ram[1891]= 7'h0;
// assign r_ram[1892]= 7'h0;
// assign r_ram[1893]= 7'h4;
// assign r_ram[1894]= 7'h8;
// assign r_ram[1895]= 7'h0;
// assign r_ram[1896]= 7'h0;
// assign r_ram[1897]= 7'h0;
// assign r_ram[1898]= 7'h0;
// assign r_ram[1899]= 7'h0;
// assign r_ram[1900]= 7'h0;
// assign r_ram[1901]= 7'h2;
// assign r_ram[1902]= 7'h0;
// assign r_ram[1903]= 7'h0;
// assign r_ram[1904]= 7'h0;
// assign r_ram[1905]= 7'h0;
// assign r_ram[1906]= 7'h0;
// assign r_ram[1907]= 7'h0;
// assign r_ram[1908]= 7'h0;
// assign r_ram[1909]= 7'h0;
// assign r_ram[1910]= 7'h11;
// assign r_ram[1911]= 7'h0;
// assign r_ram[1912]= 7'h0;
// assign r_ram[1913]= 7'h0;
// assign r_ram[1914]= 7'h0;
// assign r_ram[1915]= 7'h0;
// assign r_ram[1916]= 7'h0;
// assign r_ram[1917]= 7'h0;
// assign r_ram[1918]= 7'h0;
// assign r_ram[1919]= 7'h0;
// assign r_ram[1920]= 7'h0;
// assign r_ram[1921]= 7'h0;
// assign r_ram[1922]= 7'h0;
// assign r_ram[1923]= 7'h0;
// assign r_ram[1924]= 7'h0;
// assign r_ram[1925]= 7'h0;
// assign r_ram[1926]= 7'h0;
// assign r_ram[1927]= 7'h0;
// assign r_ram[1928]= 7'h0;
// assign r_ram[1929]= 7'h2;
// assign r_ram[1930]= 7'h0;
// assign r_ram[1931]= 7'h0;
// assign r_ram[1932]= 7'h0;
// assign r_ram[1933]= 7'h0;
// assign r_ram[1934]= 7'h4;
// assign r_ram[1935]= 7'h8;
// assign r_ram[1936]= 7'h0;
// assign r_ram[1937]= 7'h0;
// assign r_ram[1938]= 7'h0;
// assign r_ram[1939]= 7'h0;
// assign r_ram[1940]= 7'h0;
// assign r_ram[1941]= 7'h0;
// assign r_ram[1942]= 7'h0;
// assign r_ram[1943]= 7'h21;
// assign r_ram[1944]= 7'h0;
// assign r_ram[1945]= 7'h0;
// assign r_ram[1946]= 7'h0;
// assign r_ram[1947]= 7'h0;
// assign r_ram[1948]= 7'h0;
// assign r_ram[1949]= 7'h0;
// assign r_ram[1950]= 7'h0;
// assign r_ram[1951]= 7'h0;
// assign r_ram[1952]= 7'h0;
// assign r_ram[1953]= 7'h0;
// assign r_ram[1954]= 7'h0;
// assign r_ram[1955]= 7'h0;
// assign r_ram[1956]= 7'h0;
// assign r_ram[1957]= 7'h0;
// assign r_ram[1958]= 7'h0;
// assign r_ram[1959]= 7'h2;
// assign r_ram[1960]= 7'h0;
// assign r_ram[1961]= 7'h0;
// assign r_ram[1962]= 7'h0;
// assign r_ram[1963]= 7'h0;
// assign r_ram[1964]= 7'h0;
// assign r_ram[1965]= 7'h0;
// assign r_ram[1966]= 7'h0;
// assign r_ram[1967]= 7'h0;
// assign r_ram[1968]= 7'h4;
// assign r_ram[1969]= 7'h0;
// assign r_ram[1970]= 7'h0;
// assign r_ram[1971]= 7'h0;
// assign r_ram[1972]= 7'h49;
// assign r_ram[1973]= 7'h0;
// assign r_ram[1974]= 7'h0;
// assign r_ram[1975]= 7'h0;
// assign r_ram[1976]= 7'h0;
// assign r_ram[1977]= 7'h0;
// assign r_ram[1978]= 7'h0;
// assign r_ram[1979]= 7'h0;
// assign r_ram[1980]= 7'h0;
// assign r_ram[1981]= 7'h4;
// assign r_ram[1982]= 7'h8;
// assign r_ram[1983]= 7'h0;
// assign r_ram[1984]= 7'h0;
// assign r_ram[1985]= 7'h0;
// assign r_ram[1986]= 7'h0;
// assign r_ram[1987]= 7'h0;
// assign r_ram[1988]= 7'h0;
// assign r_ram[1989]= 7'h0;
// assign r_ram[1990]= 7'h0;
// assign r_ram[1991]= 7'h2;
// assign r_ram[1992]= 7'h0;
// assign r_ram[1993]= 7'h0;
// assign r_ram[1994]= 7'h0;
// assign r_ram[1995]= 7'h0;
// assign r_ram[1996]= 7'h0;
// assign r_ram[1997]= 7'h0;
// assign r_ram[1998]= 7'h0;
// assign r_ram[1999]= 7'h11;
// assign r_ram[2000]= 7'h0;
// assign r_ram[2001]= 7'h0;
// assign r_ram[2002]= 7'h0;
// assign r_ram[2003]= 7'h0;
// assign r_ram[2004]= 7'h0;
// assign r_ram[2005]= 7'h0;
// assign r_ram[2006]= 7'h0;
// assign r_ram[2007]= 7'h0;
// assign r_ram[2008]= 7'h0;
// assign r_ram[2009]= 7'h0;
// assign r_ram[2010]= 7'h0;
// assign r_ram[2011]= 7'h0;
// assign r_ram[2012]= 7'h0;
// assign r_ram[2013]= 7'h0;
// assign r_ram[2014]= 7'h0;
// assign r_ram[2015]= 7'h0;
// assign r_ram[2016]= 7'h0;
// assign r_ram[2017]= 7'h0;
// assign r_ram[2018]= 7'h2;
// assign r_ram[2019]= 7'h0;
// assign r_ram[2020]= 7'h0;
// assign r_ram[2021]= 7'h0;
// assign r_ram[2022]= 7'h0;
// assign r_ram[2023]= 7'h0;
// assign r_ram[2024]= 7'h0;
// assign r_ram[2025]= 7'h0;
// assign r_ram[2026]= 7'h0;
// assign r_ram[2027]= 7'h8;
// assign r_ram[2028]= 7'h4;
// assign r_ram[2029]= 7'h0;
// assign r_ram[2030]= 7'h0;
// assign r_ram[2031]= 7'h0;
// assign r_ram[2032]= 7'h0;
// assign r_ram[2033]= 7'h0;
// assign r_ram[2034]= 7'h21;
// assign r_ram[2035]= 7'h0;
// assign r_ram[2036]= 7'h0;
// assign r_ram[2037]= 7'h0;
// assign r_ram[2038]= 7'h0;
// assign r_ram[2039]= 7'h0;
// assign r_ram[2040]= 7'h0;
// assign r_ram[2041]= 7'h0;
// assign r_ram[2042]= 7'h0;
// assign r_ram[2043]= 7'h0;
// assign r_ram[2044]= 7'h0;
// assign r_ram[2045]= 7'h0;
// assign r_ram[2046]= 7'h0;
// assign r_ram[2047]= 7'h0;
// assign r_ram[2048]= 7'h0;
// assign r_ram[2049]= 7'h2;
// assign r_ram[2050]= 7'h0;
// assign r_ram[2051]= 7'h0;
// assign r_ram[2052]= 7'h0;
// assign r_ram[2053]= 7'h0;
// assign r_ram[2054]= 7'h0;
// assign r_ram[2055]= 7'h0;
// assign r_ram[2056]= 7'h0;
// assign r_ram[2057]= 7'h0;
// assign r_ram[2058]= 7'h0;
// assign r_ram[2059]= 7'h0;
// assign r_ram[2060]= 7'h0;
// assign r_ram[2061]= 7'h0;
// assign r_ram[2062]= 7'h8;
// assign r_ram[2063]= 7'h0;
// assign r_ram[2064]= 7'h0;
// assign r_ram[2065]= 7'h0;
// assign r_ram[2066]= 7'h4;
// assign r_ram[2067]= 7'h0;
// assign r_ram[2068]= 7'h41;
// assign r_ram[2069]= 7'h0;
// assign r_ram[2070]= 7'h0;
// assign r_ram[2071]= 7'h0;
// assign r_ram[2072]= 7'h0;
// assign r_ram[2073]= 7'h0;
// assign r_ram[2074]= 7'h4;
// assign r_ram[2075]= 7'h0;
// assign r_ram[2076]= 7'h8;
// assign r_ram[2077]= 7'h0;
// assign r_ram[2078]= 7'h0;
// assign r_ram[2079]= 7'h0;
// assign r_ram[2080]= 7'h2;
// assign r_ram[2081]= 7'h0;
// assign r_ram[2082]= 7'h0;
// assign r_ram[2083]= 7'h0;
// assign r_ram[2084]= 7'h0;
// assign r_ram[2085]= 7'h0;
// assign r_ram[2086]= 7'h0;
// assign r_ram[2087]= 7'h0;
// assign r_ram[2088]= 7'h0;
// assign r_ram[2089]= 7'h0;
// assign r_ram[2090]= 7'h11;
// assign r_ram[2091]= 7'h0;
// assign r_ram[2092]= 7'h0;
// assign r_ram[2093]= 7'h0;
// assign r_ram[2094]= 7'h0;
// assign r_ram[2095]= 7'h0;
// assign r_ram[2096]= 7'h0;
// assign r_ram[2097]= 7'h0;
// assign r_ram[2098]= 7'h0;
// assign r_ram[2099]= 7'h0;
// assign r_ram[2100]= 7'h0;
// assign r_ram[2101]= 7'h0;
// assign r_ram[2102]= 7'h0;
// assign r_ram[2103]= 7'h0;
// assign r_ram[2104]= 7'h0;
// assign r_ram[2105]= 7'h0;
// assign r_ram[2106]= 7'h0;
// assign r_ram[2107]= 7'h0;
// assign r_ram[2108]= 7'h0;
// assign r_ram[2109]= 7'h2;
// assign r_ram[2110]= 7'h0;
// assign r_ram[2111]= 7'h0;
// assign r_ram[2112]= 7'h0;
// assign r_ram[2113]= 7'h8;
// assign r_ram[2114]= 7'h0;
// assign r_ram[2115]= 7'h0;
// assign r_ram[2116]= 7'h0;
// assign r_ram[2117]= 7'h4;
// assign r_ram[2118]= 7'h0;
// assign r_ram[2119]= 7'h0;
// assign r_ram[2120]= 7'h0;
// assign r_ram[2121]= 7'h0;
// assign r_ram[2122]= 7'h0;
// assign r_ram[2123]= 7'h21;
// assign r_ram[2124]= 7'h0;
// assign r_ram[2125]= 7'h0;
// assign r_ram[2126]= 7'h0;
// assign r_ram[2127]= 7'h0;
// assign r_ram[2128]= 7'h0;
// assign r_ram[2129]= 7'h0;
// assign r_ram[2130]= 7'h0;
// assign r_ram[2131]= 7'h0;
// assign r_ram[2132]= 7'h0;
// assign r_ram[2133]= 7'h0;
// assign r_ram[2134]= 7'h0;
// assign r_ram[2135]= 7'h0;
// assign r_ram[2136]= 7'h0;
// assign r_ram[2137]= 7'h0;
// assign r_ram[2138]= 7'h0;
// assign r_ram[2139]= 7'h2;
// assign r_ram[2140]= 7'h0;
// assign r_ram[2141]= 7'h0;
// assign r_ram[2142]= 7'h0;
// assign r_ram[2143]= 7'h0;
// assign r_ram[2144]= 7'h0;
// assign r_ram[2145]= 7'h0;
// assign r_ram[2146]= 7'h0;
// assign r_ram[2147]= 7'h0;
// assign r_ram[2148]= 7'h4;
// assign r_ram[2149]= 7'h0;
// assign r_ram[2150]= 7'h8;
// assign r_ram[2151]= 7'h0;
// assign r_ram[2152]= 7'h0;
// assign r_ram[2153]= 7'h0;
// assign r_ram[2154]= 7'h41;
// assign r_ram[2155]= 7'h0;
// assign r_ram[2156]= 7'h0;
// assign r_ram[2157]= 7'h0;
// assign r_ram[2158]= 7'h0;
// assign r_ram[2159]= 7'h0;
// assign r_ram[2160]= 7'h0;
// assign r_ram[2161]= 7'h0;
// assign r_ram[2162]= 7'h8;
// assign r_ram[2163]= 7'h0;
// assign r_ram[2164]= 7'h0;
// assign r_ram[2165]= 7'h4;
// assign r_ram[2166]= 7'h0;
// assign r_ram[2167]= 7'h0;
// assign r_ram[2168]= 7'h0;
// assign r_ram[2169]= 7'h0;
// assign r_ram[2170]= 7'h2;
// assign r_ram[2171]= 7'h0;
// assign r_ram[2172]= 7'h0;
// assign r_ram[2173]= 7'h0;
// assign r_ram[2174]= 7'h0;
// assign r_ram[2175]= 7'h0;
// assign r_ram[2176]= 7'h0;
// assign r_ram[2177]= 7'h0;
// assign r_ram[2178]= 7'h0;
// assign r_ram[2179]= 7'h11;
// assign r_ram[2180]= 7'h0;
// assign r_ram[2181]= 7'h0;
// assign r_ram[2182]= 7'h0;
// assign r_ram[2183]= 7'h0;
// assign r_ram[2184]= 7'h0;
// assign r_ram[2185]= 7'h0;
// assign r_ram[2186]= 7'h0;
// assign r_ram[2187]= 7'h0;
// assign r_ram[2188]= 7'h0;
// assign r_ram[2189]= 7'h0;
// assign r_ram[2190]= 7'h0;
// assign r_ram[2191]= 7'h0;
// assign r_ram[2192]= 7'h0;
// assign r_ram[2193]= 7'h0;
// assign r_ram[2194]= 7'h0;
// assign r_ram[2195]= 7'h0;
// assign r_ram[2196]= 7'h0;
// assign r_ram[2197]= 7'h0;
// assign r_ram[2198]= 7'h0;
// assign r_ram[2199]= 7'h2;
// assign r_ram[2200]= 7'h0;
// assign r_ram[2201]= 7'h0;
// assign r_ram[2202]= 7'h0;
// assign r_ram[2203]= 7'h0;
// assign r_ram[2204]= 7'h0;
// assign r_ram[2205]= 7'h8;
// assign r_ram[2206]= 7'h4;
// assign r_ram[2207]= 7'h0;
// assign r_ram[2208]= 7'h0;
// assign r_ram[2209]= 7'h0;
// assign r_ram[2210]= 7'h0;
// assign r_ram[2211]= 7'h0;
// assign r_ram[2212]= 7'h0;
// assign r_ram[2213]= 7'h0;
// assign r_ram[2214]= 7'h21;
// assign r_ram[2215]= 7'h0;
// assign r_ram[2216]= 7'h0;
// assign r_ram[2217]= 7'h0;
// assign r_ram[2218]= 7'h0;
// assign r_ram[2219]= 7'h0;
// assign r_ram[2220]= 7'h0;
// assign r_ram[2221]= 7'h0;
// assign r_ram[2222]= 7'h0;
// assign r_ram[2223]= 7'h0;
// assign r_ram[2224]= 7'h0;
// assign r_ram[2225]= 7'h0;
// assign r_ram[2226]= 7'h0;
// assign r_ram[2227]= 7'h0;
// assign r_ram[2228]= 7'h0;
// assign r_ram[2229]= 7'h0;
// assign r_ram[2230]= 7'h2;
// assign r_ram[2231]= 7'h0;
// assign r_ram[2232]= 7'h0;
// assign r_ram[2233]= 7'h0;
// assign r_ram[2234]= 7'h0;
// assign r_ram[2235]= 7'h0;
// assign r_ram[2236]= 7'h0;
// assign r_ram[2237]= 7'h0;
// assign r_ram[2238]= 7'h0;
// assign r_ram[2239]= 7'h0;
// assign r_ram[2240]= 7'h0;
// assign r_ram[2241]= 7'h0;
// assign r_ram[2242]= 7'h4;
// assign r_ram[2243]= 7'h8;
// assign r_ram[2244]= 7'h0;
// assign r_ram[2245]= 7'h41;
// assign r_ram[2246]= 7'h0;
// assign r_ram[2247]= 7'h0;
// assign r_ram[2248]= 7'h0;
// assign r_ram[2249]= 7'h0;
assign r_ram[0]= 7'h0;
assign r_ram[1]= 7'h0;
assign r_ram[2]= 7'h0;
assign r_ram[3]= 7'h0;
assign r_ram[4]= 7'h0;
assign r_ram[5]= 7'h4;
assign r_ram[6]= 7'h8;
assign r_ram[7]= 7'h0;
assign r_ram[8]= 7'h0;
assign r_ram[9]= 7'h0;
assign r_ram[10]= 7'h0;
assign r_ram[11]= 7'h2;
assign r_ram[12]= 7'h0;
assign r_ram[13]= 7'h0;
assign r_ram[14]= 7'h0;
assign r_ram[15]= 7'h0;
assign r_ram[16]= 7'h0;
assign r_ram[17]= 7'h0;
assign r_ram[18]= 7'h0;
assign r_ram[19]= 7'h0;
assign r_ram[20]= 7'h0;
assign r_ram[21]= 7'h0;
assign r_ram[22]= 7'h0;
assign r_ram[23]= 7'h11;
assign r_ram[24]= 7'h0;
assign r_ram[25]= 7'h0;
assign r_ram[26]= 7'h0;
assign r_ram[27]= 7'h0;
assign r_ram[28]= 7'h0;
assign r_ram[29]= 7'h0;
assign r_ram[30]= 7'h0;
assign r_ram[31]= 7'h0;
assign r_ram[32]= 7'h0;
assign r_ram[33]= 7'h0;
assign r_ram[34]= 7'h0;
assign r_ram[35]= 7'h0;
assign r_ram[36]= 7'h0;
assign r_ram[37]= 7'h0;
assign r_ram[38]= 7'h0;
assign r_ram[39]= 7'h0;
assign r_ram[40]= 7'h0;
assign r_ram[41]= 7'h2;
assign r_ram[42]= 7'h0;
assign r_ram[43]= 7'h0;
assign r_ram[44]= 7'h0;
assign r_ram[45]= 7'h0;
assign r_ram[46]= 7'h0;
assign r_ram[47]= 7'h0;
assign r_ram[48]= 7'hc;
assign r_ram[49]= 7'h0;
assign r_ram[50]= 7'h0;
assign r_ram[51]= 7'h0;
assign r_ram[52]= 7'h0;
assign r_ram[53]= 7'h0;
assign r_ram[54]= 7'h0;
assign r_ram[55]= 7'h0;
assign r_ram[56]= 7'h0;
assign r_ram[57]= 7'h21;
assign r_ram[58]= 7'h0;
assign r_ram[59]= 7'h0;
assign r_ram[60]= 7'h0;
assign r_ram[61]= 7'h0;
assign r_ram[62]= 7'h0;
assign r_ram[63]= 7'h0;
assign r_ram[64]= 7'h0;
assign r_ram[65]= 7'h0;
assign r_ram[66]= 7'h0;
assign r_ram[67]= 7'h0;
assign r_ram[68]= 7'h0;
assign r_ram[69]= 7'h0;
assign r_ram[70]= 7'h0;
assign r_ram[71]= 7'h2;
assign r_ram[72]= 7'h0;
assign r_ram[73]= 7'h0;
assign r_ram[74]= 7'h0;
assign r_ram[75]= 7'h0;
assign r_ram[76]= 7'h0;
assign r_ram[77]= 7'h0;
assign r_ram[78]= 7'h0;
assign r_ram[79]= 7'h0;
assign r_ram[80]= 7'h0;
assign r_ram[81]= 7'h0;
assign r_ram[82]= 7'h0;
assign r_ram[83]= 7'h4;
assign r_ram[84]= 7'h0;
assign r_ram[85]= 7'h0;
assign r_ram[86]= 7'h1;
assign r_ram[87]= 7'h0;
assign r_ram[88]= 7'h0;
assign r_ram[89]= 7'h48;
assign r_ram[90]= 7'h0;
assign r_ram[91]= 7'h0;
assign r_ram[92]= 7'h0;
assign r_ram[93]= 7'h0;
assign r_ram[94]= 7'h0;
assign r_ram[95]= 7'h4;
assign r_ram[96]= 7'h8;
assign r_ram[97]= 7'h0;
assign r_ram[98]= 7'h0;
assign r_ram[99]= 7'h0;
assign r_ram[100]= 7'h2;
assign r_ram[101]= 7'h0;
assign r_ram[102]= 7'h0;
assign r_ram[103]= 7'h0;
assign r_ram[104]= 7'h0;
assign r_ram[105]= 7'h0;
assign r_ram[106]= 7'h0;
assign r_ram[107]= 7'h0;
assign r_ram[108]= 7'h0;
assign r_ram[109]= 7'h0;
assign r_ram[110]= 7'h0;
assign r_ram[111]= 7'h0;
assign r_ram[112]= 7'h0;
assign r_ram[113]= 7'h11;
assign r_ram[114]= 7'h0;
assign r_ram[115]= 7'h0;
assign r_ram[116]= 7'h0;
assign r_ram[117]= 7'h0;
assign r_ram[118]= 7'h0;
assign r_ram[119]= 7'h0;
assign r_ram[120]= 7'h0;
assign r_ram[121]= 7'h0;
assign r_ram[122]= 7'h0;
assign r_ram[123]= 7'h0;
assign r_ram[124]= 7'h0;
assign r_ram[125]= 7'h0;
assign r_ram[126]= 7'h0;
assign r_ram[127]= 7'h0;
assign r_ram[128]= 7'h0;
assign r_ram[129]= 7'h0;
assign r_ram[130]= 7'h0;
assign r_ram[131]= 7'h2;
assign r_ram[132]= 7'h0;
assign r_ram[133]= 7'h0;
assign r_ram[134]= 7'h0;
assign r_ram[135]= 7'h0;
assign r_ram[136]= 7'h0;
assign r_ram[137]= 7'h4;
assign r_ram[138]= 7'h0;
assign r_ram[139]= 7'h8;
assign r_ram[140]= 7'h0;
assign r_ram[141]= 7'h0;
assign r_ram[142]= 7'h0;
assign r_ram[143]= 7'h0;
assign r_ram[144]= 7'h0;
assign r_ram[145]= 7'h0;
assign r_ram[146]= 7'h21;
assign r_ram[147]= 7'h0;
assign r_ram[148]= 7'h0;
assign r_ram[149]= 7'h0;
assign r_ram[150]= 7'h0;
assign r_ram[151]= 7'h0;
assign r_ram[152]= 7'h0;
assign r_ram[153]= 7'h0;
assign r_ram[154]= 7'h0;
assign r_ram[155]= 7'h0;
assign r_ram[156]= 7'h0;
assign r_ram[157]= 7'h0;
assign r_ram[158]= 7'h0;
assign r_ram[159]= 7'h0;
assign r_ram[160]= 7'h2;
assign r_ram[161]= 7'h0;
assign r_ram[162]= 7'h0;
assign r_ram[163]= 7'h0;
assign r_ram[164]= 7'h0;
assign r_ram[165]= 7'h0;
assign r_ram[166]= 7'h0;
assign r_ram[167]= 7'h0;
assign r_ram[168]= 7'h0;
assign r_ram[169]= 7'h4;
assign r_ram[170]= 7'h0;
assign r_ram[171]= 7'h0;
assign r_ram[172]= 7'h0;
assign r_ram[173]= 7'h8;
assign r_ram[174]= 7'h0;
assign r_ram[175]= 7'h41;
assign r_ram[176]= 7'h0;
assign r_ram[177]= 7'h0;
assign r_ram[178]= 7'h0;
assign r_ram[179]= 7'h0;
assign r_ram[180]= 7'h0;
assign r_ram[181]= 7'h0;
assign r_ram[182]= 7'h0;
assign r_ram[183]= 7'h0;
assign r_ram[184]= 7'h0;
assign r_ram[185]= 7'h4;
assign r_ram[186]= 7'h8;
assign r_ram[187]= 7'h0;
assign r_ram[188]= 7'h0;
assign r_ram[189]= 7'h0;
assign r_ram[190]= 7'h0;
assign r_ram[191]= 7'h2;
assign r_ram[192]= 7'h0;
assign r_ram[193]= 7'h0;
assign r_ram[194]= 7'h0;
assign r_ram[195]= 7'h0;
assign r_ram[196]= 7'h0;
assign r_ram[197]= 7'h0;
assign r_ram[198]= 7'h0;
assign r_ram[199]= 7'h0;
assign r_ram[200]= 7'h0;
assign r_ram[201]= 7'h0;
assign r_ram[202]= 7'h0;
assign r_ram[203]= 7'h11;
assign r_ram[204]= 7'h0;
assign r_ram[205]= 7'h0;
assign r_ram[206]= 7'h0;
assign r_ram[207]= 7'h0;
assign r_ram[208]= 7'h0;
assign r_ram[209]= 7'h0;
assign r_ram[210]= 7'h0;
assign r_ram[211]= 7'h0;
assign r_ram[212]= 7'h0;
assign r_ram[213]= 7'h0;
assign r_ram[214]= 7'h0;
assign r_ram[215]= 7'h0;
assign r_ram[216]= 7'h0;
assign r_ram[217]= 7'h0;
assign r_ram[218]= 7'h0;
assign r_ram[219]= 7'h0;
assign r_ram[220]= 7'h2;
assign r_ram[221]= 7'h0;
assign r_ram[222]= 7'h0;
assign r_ram[223]= 7'h0;
assign r_ram[224]= 7'h0;
assign r_ram[225]= 7'h0;
assign r_ram[226]= 7'h0;
assign r_ram[227]= 7'h0;
assign r_ram[228]= 7'h0;
assign r_ram[229]= 7'hc;
assign r_ram[230]= 7'h0;
assign r_ram[231]= 7'h0;
assign r_ram[232]= 7'h0;
assign r_ram[233]= 7'h0;
assign r_ram[234]= 7'h0;
assign r_ram[235]= 7'h0;
assign r_ram[236]= 7'h0;
assign r_ram[237]= 7'h21;
assign r_ram[238]= 7'h0;
assign r_ram[239]= 7'h0;
assign r_ram[240]= 7'h0;
assign r_ram[241]= 7'h0;
assign r_ram[242]= 7'h0;
assign r_ram[243]= 7'h0;
assign r_ram[244]= 7'h0;
assign r_ram[245]= 7'h0;
assign r_ram[246]= 7'h0;
assign r_ram[247]= 7'h0;
assign r_ram[248]= 7'h0;
assign r_ram[249]= 7'h0;
assign r_ram[250]= 7'h2;
assign r_ram[251]= 7'h0;
assign r_ram[252]= 7'h0;
assign r_ram[253]= 7'h0;
assign r_ram[254]= 7'h0;
assign r_ram[255]= 7'h0;
assign r_ram[256]= 7'h0;
assign r_ram[257]= 7'h0;
assign r_ram[258]= 7'h0;
assign r_ram[259]= 7'h0;
assign r_ram[260]= 7'h0;
assign r_ram[261]= 7'h0;
assign r_ram[262]= 7'h4;
assign r_ram[263]= 7'h0;
assign r_ram[264]= 7'h0;
assign r_ram[265]= 7'h8;
assign r_ram[266]= 7'h0;
assign r_ram[267]= 7'h41;
assign r_ram[268]= 7'h0;
assign r_ram[269]= 7'h0;
assign r_ram[270]= 7'h0;
assign r_ram[271]= 7'h0;
assign r_ram[272]= 7'h0;
assign r_ram[273]= 7'h0;
assign r_ram[274]= 7'h0;
assign r_ram[275]= 7'h0;
assign r_ram[276]= 7'hc;
assign r_ram[277]= 7'h0;
assign r_ram[278]= 7'h0;
assign r_ram[279]= 7'h0;
assign r_ram[280]= 7'h2;
assign r_ram[281]= 7'h0;
assign r_ram[282]= 7'h0;
assign r_ram[283]= 7'h0;
assign r_ram[284]= 7'h0;
assign r_ram[285]= 7'h0;
assign r_ram[286]= 7'h0;
assign r_ram[287]= 7'h0;
assign r_ram[288]= 7'h0;
assign r_ram[289]= 7'h0;
assign r_ram[290]= 7'h0;
assign r_ram[291]= 7'h0;
assign r_ram[292]= 7'h11;
assign r_ram[293]= 7'h0;
assign r_ram[294]= 7'h0;
assign r_ram[295]= 7'h0;
assign r_ram[296]= 7'h0;
assign r_ram[297]= 7'h0;
assign r_ram[298]= 7'h0;
assign r_ram[299]= 7'h0;
assign r_ram[300]= 7'h0;
assign r_ram[301]= 7'h0;
assign r_ram[302]= 7'h0;
assign r_ram[303]= 7'h0;
assign r_ram[304]= 7'h0;
assign r_ram[305]= 7'h0;
assign r_ram[306]= 7'h0;
assign r_ram[307]= 7'h0;
assign r_ram[308]= 7'h0;
assign r_ram[309]= 7'h2;
assign r_ram[310]= 7'h0;
assign r_ram[311]= 7'h0;
assign r_ram[312]= 7'h0;
assign r_ram[313]= 7'h0;
assign r_ram[314]= 7'h0;
assign r_ram[315]= 7'h4;
assign r_ram[316]= 7'h0;
assign r_ram[317]= 7'h8;
assign r_ram[318]= 7'h0;
assign r_ram[319]= 7'h0;
assign r_ram[320]= 7'h0;
assign r_ram[321]= 7'h0;
assign r_ram[322]= 7'h0;
assign r_ram[323]= 7'h0;
assign r_ram[324]= 7'h21;
assign r_ram[325]= 7'h0;
assign r_ram[326]= 7'h0;
assign r_ram[327]= 7'h0;
assign r_ram[328]= 7'h0;
assign r_ram[329]= 7'h0;
assign r_ram[330]= 7'h0;
assign r_ram[331]= 7'h0;
assign r_ram[332]= 7'h0;
assign r_ram[333]= 7'h0;
assign r_ram[334]= 7'h0;
assign r_ram[335]= 7'h0;
assign r_ram[336]= 7'h0;
assign r_ram[337]= 7'h0;
assign r_ram[338]= 7'h0;
assign r_ram[339]= 7'h0;
assign r_ram[340]= 7'h2;
assign r_ram[341]= 7'h0;
assign r_ram[342]= 7'h0;
assign r_ram[343]= 7'h0;
assign r_ram[344]= 7'h0;
assign r_ram[345]= 7'h0;
assign r_ram[346]= 7'h0;
assign r_ram[347]= 7'h0;
assign r_ram[348]= 7'h0;
assign r_ram[349]= 7'h0;
assign r_ram[350]= 7'h0;
assign r_ram[351]= 7'h4;
assign r_ram[352]= 7'h8;
assign r_ram[353]= 7'h0;
assign r_ram[354]= 7'h0;
assign r_ram[355]= 7'h0;
assign r_ram[356]= 7'h41;
assign r_ram[357]= 7'h0;
assign r_ram[358]= 7'h0;
assign r_ram[359]= 7'h0;
assign r_ram[360]= 7'h0;
assign r_ram[361]= 7'h0;
assign r_ram[362]= 7'h0;
assign r_ram[363]= 7'h0;
assign r_ram[364]= 7'h0;
assign r_ram[365]= 7'h4;
assign r_ram[366]= 7'h8;
assign r_ram[367]= 7'h0;
assign r_ram[368]= 7'h0;
assign r_ram[369]= 7'h0;
assign r_ram[370]= 7'h0;
assign r_ram[371]= 7'h2;
assign r_ram[372]= 7'h0;
assign r_ram[373]= 7'h0;
assign r_ram[374]= 7'h0;
assign r_ram[375]= 7'h0;
assign r_ram[376]= 7'h0;
assign r_ram[377]= 7'h0;
assign r_ram[378]= 7'h0;
assign r_ram[379]= 7'h0;
assign r_ram[380]= 7'h0;
assign r_ram[381]= 7'h0;
assign r_ram[382]= 7'h0;
assign r_ram[383]= 7'h11;
assign r_ram[384]= 7'h0;
assign r_ram[385]= 7'h0;
assign r_ram[386]= 7'h0;
assign r_ram[387]= 7'h0;
assign r_ram[388]= 7'h0;
assign r_ram[389]= 7'h0;
assign r_ram[390]= 7'h0;
assign r_ram[391]= 7'h0;
assign r_ram[392]= 7'h0;
assign r_ram[393]= 7'h0;
assign r_ram[394]= 7'h0;
assign r_ram[395]= 7'h0;
assign r_ram[396]= 7'h0;
assign r_ram[397]= 7'h0;
assign r_ram[398]= 7'h0;
assign r_ram[399]= 7'h0;
assign r_ram[400]= 7'h2;
assign r_ram[401]= 7'h0;
assign r_ram[402]= 7'h0;
assign r_ram[403]= 7'h0;
assign r_ram[404]= 7'h0;
assign r_ram[405]= 7'h0;
assign r_ram[406]= 7'h0;
assign r_ram[407]= 7'h4;
assign r_ram[408]= 7'h0;
assign r_ram[409]= 7'h8;
assign r_ram[410]= 7'h0;
assign r_ram[411]= 7'h0;
assign r_ram[412]= 7'h0;
assign r_ram[413]= 7'h0;
assign r_ram[414]= 7'h0;
assign r_ram[415]= 7'h0;
assign r_ram[416]= 7'h21;
assign r_ram[417]= 7'h0;
assign r_ram[418]= 7'h0;
assign r_ram[419]= 7'h0;
assign r_ram[420]= 7'h0;
assign r_ram[421]= 7'h0;
assign r_ram[422]= 7'h0;
assign r_ram[423]= 7'h0;
assign r_ram[424]= 7'h0;
assign r_ram[425]= 7'h0;
assign r_ram[426]= 7'h0;
assign r_ram[427]= 7'h0;
assign r_ram[428]= 7'h0;
assign r_ram[429]= 7'h0;
assign r_ram[430]= 7'h2;
assign r_ram[431]= 7'h0;
assign r_ram[432]= 7'h0;
assign r_ram[433]= 7'h0;
assign r_ram[434]= 7'h0;
assign r_ram[435]= 7'h0;
assign r_ram[436]= 7'h0;
assign r_ram[437]= 7'h0;
assign r_ram[438]= 7'h0;
assign r_ram[439]= 7'h0;
assign r_ram[440]= 7'h0;
assign r_ram[441]= 7'h0;
assign r_ram[442]= 7'h4;
assign r_ram[443]= 7'h0;
assign r_ram[444]= 7'h0;
assign r_ram[445]= 7'h0;
assign r_ram[446]= 7'h49;
assign r_ram[447]= 7'h0;
assign r_ram[448]= 7'h0;
assign r_ram[449]= 7'h0;
assign r_ram[450]= 7'h0;
assign r_ram[451]= 7'h0;
assign r_ram[452]= 7'h0;
assign r_ram[453]= 7'h0;
assign r_ram[454]= 7'h0;
assign r_ram[455]= 7'h0;
assign r_ram[456]= 7'h4;
assign r_ram[457]= 7'h0;
assign r_ram[458]= 7'h8;
assign r_ram[459]= 7'h0;
assign r_ram[460]= 7'h0;
assign r_ram[461]= 7'h2;
assign r_ram[462]= 7'h0;
assign r_ram[463]= 7'h0;
assign r_ram[464]= 7'h0;
assign r_ram[465]= 7'h0;
assign r_ram[466]= 7'h0;
assign r_ram[467]= 7'h0;
assign r_ram[468]= 7'h0;
assign r_ram[469]= 7'h0;
assign r_ram[470]= 7'h0;
assign r_ram[471]= 7'h0;
assign r_ram[472]= 7'h0;
assign r_ram[473]= 7'h0;
assign r_ram[474]= 7'h11;
assign r_ram[475]= 7'h0;
assign r_ram[476]= 7'h0;
assign r_ram[477]= 7'h0;
assign r_ram[478]= 7'h0;
assign r_ram[479]= 7'h0;
assign r_ram[480]= 7'h0;
assign r_ram[481]= 7'h0;
assign r_ram[482]= 7'h0;
assign r_ram[483]= 7'h0;
assign r_ram[484]= 7'h0;
assign r_ram[485]= 7'h0;
assign r_ram[486]= 7'h0;
assign r_ram[487]= 7'h0;
assign r_ram[488]= 7'h0;
assign r_ram[489]= 7'h0;
assign r_ram[490]= 7'h2;
assign r_ram[491]= 7'h0;
assign r_ram[492]= 7'h0;
assign r_ram[493]= 7'h0;
assign r_ram[494]= 7'h0;
assign r_ram[495]= 7'h0;
assign r_ram[496]= 7'h0;
assign r_ram[497]= 7'hc;
assign r_ram[498]= 7'h0;
assign r_ram[499]= 7'h0;
assign r_ram[500]= 7'h0;
assign r_ram[501]= 7'h0;
assign r_ram[502]= 7'h0;
assign r_ram[503]= 7'h0;
assign r_ram[504]= 7'h0;
assign r_ram[505]= 7'h21;
assign r_ram[506]= 7'h0;
assign r_ram[507]= 7'h0;
assign r_ram[508]= 7'h0;
assign r_ram[509]= 7'h0;
assign r_ram[510]= 7'h0;
assign r_ram[511]= 7'h0;
assign r_ram[512]= 7'h0;
assign r_ram[513]= 7'h0;
assign r_ram[514]= 7'h0;
assign r_ram[515]= 7'h0;
assign r_ram[516]= 7'h0;
assign r_ram[517]= 7'h0;
assign r_ram[518]= 7'h0;
assign r_ram[519]= 7'h0;
assign r_ram[520]= 7'h2;
assign r_ram[521]= 7'h0;
assign r_ram[522]= 7'h0;
assign r_ram[523]= 7'h0;
assign r_ram[524]= 7'h0;
assign r_ram[525]= 7'h0;
assign r_ram[526]= 7'h0;
assign r_ram[527]= 7'h0;
assign r_ram[528]= 7'h0;
assign r_ram[529]= 7'h0;
assign r_ram[530]= 7'h0;
assign r_ram[531]= 7'h0;
assign r_ram[532]= 7'h0;
assign r_ram[533]= 7'h0;
assign r_ram[534]= 7'h0;
assign r_ram[535]= 7'hc;
assign r_ram[536]= 7'h0;
assign r_ram[537]= 7'h0;
assign r_ram[538]= 7'h41;
assign r_ram[539]= 7'h0;
assign r_ram[540]= 7'h0;
assign r_ram[541]= 7'h0;
assign r_ram[542]= 7'h0;
assign r_ram[543]= 7'h0;
assign r_ram[544]= 7'h0;
assign r_ram[545]= 7'h4;
assign r_ram[546]= 7'h0;
assign r_ram[547]= 7'h8;
assign r_ram[548]= 7'h0;
assign r_ram[549]= 7'h0;
assign r_ram[550]= 7'h0;
assign r_ram[551]= 7'h2;
assign r_ram[552]= 7'h0;
assign r_ram[553]= 7'h0;
assign r_ram[554]= 7'h0;
assign r_ram[555]= 7'h0;
assign r_ram[556]= 7'h0;
assign r_ram[557]= 7'h0;
assign r_ram[558]= 7'h0;
assign r_ram[559]= 7'h0;
assign r_ram[560]= 7'h0;
assign r_ram[561]= 7'h0;
assign r_ram[562]= 7'h11;
assign r_ram[563]= 7'h0;
assign r_ram[564]= 7'h0;
assign r_ram[565]= 7'h0;
assign r_ram[566]= 7'h0;
assign r_ram[567]= 7'h0;
assign r_ram[568]= 7'h0;
assign r_ram[569]= 7'h0;
assign r_ram[570]= 7'h0;
assign r_ram[571]= 7'h0;
assign r_ram[572]= 7'h0;
assign r_ram[573]= 7'h0;
assign r_ram[574]= 7'h0;
assign r_ram[575]= 7'h0;
assign r_ram[576]= 7'h0;
assign r_ram[577]= 7'h0;
assign r_ram[578]= 7'h0;
assign r_ram[579]= 7'h0;
assign r_ram[580]= 7'h0;
assign r_ram[581]= 7'h2;
assign r_ram[582]= 7'h0;
assign r_ram[583]= 7'h0;
assign r_ram[584]= 7'h0;
assign r_ram[585]= 7'h0;
assign r_ram[586]= 7'h0;
assign r_ram[587]= 7'h0;
assign r_ram[588]= 7'h4;
assign r_ram[589]= 7'h0;
assign r_ram[590]= 7'h8;
assign r_ram[591]= 7'h0;
assign r_ram[592]= 7'h0;
assign r_ram[593]= 7'h0;
assign r_ram[594]= 7'h0;
assign r_ram[595]= 7'h0;
assign r_ram[596]= 7'h21;
assign r_ram[597]= 7'h0;
assign r_ram[598]= 7'h0;
assign r_ram[599]= 7'h0;
assign r_ram[600]= 7'h0;
assign r_ram[601]= 7'h0;
assign r_ram[602]= 7'h0;
assign r_ram[603]= 7'h0;
assign r_ram[604]= 7'h0;
assign r_ram[605]= 7'h0;
assign r_ram[606]= 7'h0;
assign r_ram[607]= 7'h0;
assign r_ram[608]= 7'h0;
assign r_ram[609]= 7'h0;
assign r_ram[610]= 7'h2;
assign r_ram[611]= 7'h0;
assign r_ram[612]= 7'h0;
assign r_ram[613]= 7'h0;
assign r_ram[614]= 7'h0;
assign r_ram[615]= 7'h0;
assign r_ram[616]= 7'h0;
assign r_ram[617]= 7'h4;
assign r_ram[618]= 7'h0;
assign r_ram[619]= 7'h0;
assign r_ram[620]= 7'h0;
assign r_ram[621]= 7'h8;
assign r_ram[622]= 7'h0;
assign r_ram[623]= 7'h41;
assign r_ram[624]= 7'h0;
assign r_ram[625]= 7'h0;
assign r_ram[626]= 7'h0;
assign r_ram[627]= 7'h0;
assign r_ram[628]= 7'h0;
assign r_ram[629]= 7'h0;
assign r_ram[630]= 7'h0;
assign r_ram[631]= 7'h0;
assign r_ram[632]= 7'h0;
assign r_ram[633]= 7'h0;
assign r_ram[634]= 7'h0;
assign r_ram[635]= 7'h0;
assign r_ram[636]= 7'hc;
assign r_ram[637]= 7'h0;
assign r_ram[638]= 7'h0;
assign r_ram[639]= 7'h0;
assign r_ram[640]= 7'h0;
assign r_ram[641]= 7'h2;
assign r_ram[642]= 7'h0;
assign r_ram[643]= 7'h0;
assign r_ram[644]= 7'h0;
assign r_ram[645]= 7'h0;
assign r_ram[646]= 7'h0;
assign r_ram[647]= 7'h0;
assign r_ram[648]= 7'h0;
assign r_ram[649]= 7'h0;
assign r_ram[650]= 7'h0;
assign r_ram[651]= 7'h0;
assign r_ram[652]= 7'h0;
assign r_ram[653]= 7'h11;
assign r_ram[654]= 7'h0;
assign r_ram[655]= 7'h0;
assign r_ram[656]= 7'h0;
assign r_ram[657]= 7'h0;
assign r_ram[658]= 7'h0;
assign r_ram[659]= 7'h0;
assign r_ram[660]= 7'h0;
assign r_ram[661]= 7'h0;
assign r_ram[662]= 7'h0;
assign r_ram[663]= 7'h0;
assign r_ram[664]= 7'h0;
assign r_ram[665]= 7'h0;
assign r_ram[666]= 7'h0;
assign r_ram[667]= 7'h0;
assign r_ram[668]= 7'h0;
assign r_ram[669]= 7'h0;
assign r_ram[670]= 7'h2;
assign r_ram[671]= 7'h0;
assign r_ram[672]= 7'h4;
assign r_ram[673]= 7'h0;
assign r_ram[674]= 7'h8;
assign r_ram[675]= 7'h0;
assign r_ram[676]= 7'h0;
assign r_ram[677]= 7'h0;
assign r_ram[678]= 7'h0;
assign r_ram[679]= 7'h0;
assign r_ram[680]= 7'h0;
assign r_ram[681]= 7'h0;
assign r_ram[682]= 7'h0;
assign r_ram[683]= 7'h21;
assign r_ram[684]= 7'h0;
assign r_ram[685]= 7'h0;
assign r_ram[686]= 7'h0;
assign r_ram[687]= 7'h0;
assign r_ram[688]= 7'h0;
assign r_ram[689]= 7'h0;
assign r_ram[690]= 7'h0;
assign r_ram[691]= 7'h0;
assign r_ram[692]= 7'h0;
assign r_ram[693]= 7'h0;
assign r_ram[694]= 7'h0;
assign r_ram[695]= 7'h0;
assign r_ram[696]= 7'h0;
assign r_ram[697]= 7'h0;
assign r_ram[698]= 7'h0;
assign r_ram[699]= 7'h0;
assign r_ram[700]= 7'h2;
assign r_ram[701]= 7'h0;
assign r_ram[702]= 7'h0;
assign r_ram[703]= 7'h0;
assign r_ram[704]= 7'h0;
assign r_ram[705]= 7'h0;
assign r_ram[706]= 7'h0;
assign r_ram[707]= 7'h0;
assign r_ram[708]= 7'h0;
assign r_ram[709]= 7'h0;
assign r_ram[710]= 7'h0;
assign r_ram[711]= 7'h0;
assign r_ram[712]= 7'h8;
assign r_ram[713]= 7'h0;
assign r_ram[714]= 7'h4;
assign r_ram[715]= 7'h0;
assign r_ram[716]= 7'h0;
assign r_ram[717]= 7'h0;
assign r_ram[718]= 7'h41;
assign r_ram[719]= 7'h0;
assign r_ram[720]= 7'h0;
assign r_ram[721]= 7'h0;
assign r_ram[722]= 7'h0;
assign r_ram[723]= 7'h0;
assign r_ram[724]= 7'h0;
assign r_ram[725]= 7'h4;
assign r_ram[726]= 7'h8;
assign r_ram[727]= 7'h0;
assign r_ram[728]= 7'h0;
assign r_ram[729]= 7'h0;
assign r_ram[730]= 7'h2;
assign r_ram[731]= 7'h0;
assign r_ram[732]= 7'h0;
assign r_ram[733]= 7'h0;
assign r_ram[734]= 7'h0;
assign r_ram[735]= 7'h0;
assign r_ram[736]= 7'h0;
assign r_ram[737]= 7'h0;
assign r_ram[738]= 7'h0;
assign r_ram[739]= 7'h0;
assign r_ram[740]= 7'h0;
assign r_ram[741]= 7'h0;
assign r_ram[742]= 7'h11;
assign r_ram[743]= 7'h0;
assign r_ram[744]= 7'h0;
assign r_ram[745]= 7'h0;
assign r_ram[746]= 7'h0;
assign r_ram[747]= 7'h0;
assign r_ram[748]= 7'h0;
assign r_ram[749]= 7'h0;
assign r_ram[750]= 7'h0;
assign r_ram[751]= 7'h0;
assign r_ram[752]= 7'h0;
assign r_ram[753]= 7'h0;
assign r_ram[754]= 7'h0;
assign r_ram[755]= 7'h0;
assign r_ram[756]= 7'h0;
assign r_ram[757]= 7'h0;
assign r_ram[758]= 7'h0;
assign r_ram[759]= 7'h0;
assign r_ram[760]= 7'h2;
assign r_ram[761]= 7'h0;
assign r_ram[762]= 7'h0;
assign r_ram[763]= 7'h0;
assign r_ram[764]= 7'h0;
assign r_ram[765]= 7'h0;
assign r_ram[766]= 7'h0;
assign r_ram[767]= 7'hc;
assign r_ram[768]= 7'h0;
assign r_ram[769]= 7'h0;
assign r_ram[770]= 7'h0;
assign r_ram[771]= 7'h0;
assign r_ram[772]= 7'h0;
assign r_ram[773]= 7'h0;
assign r_ram[774]= 7'h0;
assign r_ram[775]= 7'h0;
assign r_ram[776]= 7'h21;
assign r_ram[777]= 7'h0;
assign r_ram[778]= 7'h0;
assign r_ram[779]= 7'h0;
assign r_ram[780]= 7'h0;
assign r_ram[781]= 7'h0;
assign r_ram[782]= 7'h0;
assign r_ram[783]= 7'h0;
assign r_ram[784]= 7'h0;
assign r_ram[785]= 7'h0;
assign r_ram[786]= 7'h0;
assign r_ram[787]= 7'h0;
assign r_ram[788]= 7'h0;
assign r_ram[789]= 7'h0;
assign r_ram[790]= 7'h2;
assign r_ram[791]= 7'h0;
assign r_ram[792]= 7'h0;
assign r_ram[793]= 7'h0;
assign r_ram[794]= 7'h0;
assign r_ram[795]= 7'h0;
assign r_ram[796]= 7'h0;
assign r_ram[797]= 7'h0;
assign r_ram[798]= 7'h0;
assign r_ram[799]= 7'h0;
assign r_ram[800]= 7'h0;
assign r_ram[801]= 7'h0;
assign r_ram[802]= 7'hc;
assign r_ram[803]= 7'h0;
assign r_ram[804]= 7'h0;
assign r_ram[805]= 7'h0;
assign r_ram[806]= 7'h41;
assign r_ram[807]= 7'h0;
assign r_ram[808]= 7'h0;
assign r_ram[809]= 7'h0;
assign r_ram[810]= 7'h0;
assign r_ram[811]= 7'h0;
assign r_ram[812]= 7'h0;
assign r_ram[813]= 7'h0;
assign r_ram[814]= 7'h0;
assign r_ram[815]= 7'h8;
assign r_ram[816]= 7'h4;
assign r_ram[817]= 7'h0;
assign r_ram[818]= 7'h0;
assign r_ram[819]= 7'h0;
assign r_ram[820]= 7'h2;
assign r_ram[821]= 7'h0;
assign r_ram[822]= 7'h0;
assign r_ram[823]= 7'h0;
assign r_ram[824]= 7'h0;
assign r_ram[825]= 7'h0;
assign r_ram[826]= 7'h0;
assign r_ram[827]= 7'h0;
assign r_ram[828]= 7'h0;
assign r_ram[829]= 7'h0;
assign r_ram[830]= 7'h0;
assign r_ram[831]= 7'h0;
assign r_ram[832]= 7'h0;
assign r_ram[833]= 7'h11;
assign r_ram[834]= 7'h0;
assign r_ram[835]= 7'h0;
assign r_ram[836]= 7'h0;
assign r_ram[837]= 7'h0;
assign r_ram[838]= 7'h0;
assign r_ram[839]= 7'h0;
assign r_ram[840]= 7'h0;
assign r_ram[841]= 7'h0;
assign r_ram[842]= 7'h0;
assign r_ram[843]= 7'h0;
assign r_ram[844]= 7'h0;
assign r_ram[845]= 7'h0;
assign r_ram[846]= 7'h0;
assign r_ram[847]= 7'h0;
assign r_ram[848]= 7'h0;
assign r_ram[849]= 7'h0;
assign r_ram[850]= 7'h2;
assign r_ram[851]= 7'h0;
assign r_ram[852]= 7'h0;
assign r_ram[853]= 7'h0;
assign r_ram[854]= 7'h0;
assign r_ram[855]= 7'h4;
assign r_ram[856]= 7'h0;
assign r_ram[857]= 7'h0;
assign r_ram[858]= 7'h8;
assign r_ram[859]= 7'h0;
assign r_ram[860]= 7'h0;
assign r_ram[861]= 7'h0;
assign r_ram[862]= 7'h0;
assign r_ram[863]= 7'h0;
assign r_ram[864]= 7'h21;
assign r_ram[865]= 7'h0;
assign r_ram[866]= 7'h0;
assign r_ram[867]= 7'h0;
assign r_ram[868]= 7'h0;
assign r_ram[869]= 7'h0;
assign r_ram[870]= 7'h0;
assign r_ram[871]= 7'h0;
assign r_ram[872]= 7'h0;
assign r_ram[873]= 7'h0;
assign r_ram[874]= 7'h0;
assign r_ram[875]= 7'h0;
assign r_ram[876]= 7'h0;
assign r_ram[877]= 7'h0;
assign r_ram[878]= 7'h0;
assign r_ram[879]= 7'h0;
assign r_ram[880]= 7'h0;
assign r_ram[881]= 7'h2;
assign r_ram[882]= 7'h0;
assign r_ram[883]= 7'h0;
assign r_ram[884]= 7'h0;
assign r_ram[885]= 7'h0;
assign r_ram[886]= 7'h0;
assign r_ram[887]= 7'h0;
assign r_ram[888]= 7'h0;
assign r_ram[889]= 7'h0;
assign r_ram[890]= 7'h0;
assign r_ram[891]= 7'h0;
assign r_ram[892]= 7'h0;
assign r_ram[893]= 7'h4;
assign r_ram[894]= 7'h0;
assign r_ram[895]= 7'h0;
assign r_ram[896]= 7'h0;
assign r_ram[897]= 7'h1;
assign r_ram[898]= 7'h0;
assign r_ram[899]= 7'h48;
assign r_ram[900]= 7'h0;
assign r_ram[901]= 7'h0;
assign r_ram[902]= 7'h0;
assign r_ram[903]= 7'h0;
assign r_ram[904]= 7'h0;
assign r_ram[905]= 7'h0;
assign r_ram[906]= 7'hc;
assign r_ram[907]= 7'h0;
assign r_ram[908]= 7'h0;
assign r_ram[909]= 7'h0;
assign r_ram[910]= 7'h0;
assign r_ram[911]= 7'h2;
assign r_ram[912]= 7'h0;
assign r_ram[913]= 7'h0;
assign r_ram[914]= 7'h0;
assign r_ram[915]= 7'h0;
assign r_ram[916]= 7'h0;
assign r_ram[917]= 7'h0;
assign r_ram[918]= 7'h0;
assign r_ram[919]= 7'h0;
assign r_ram[920]= 7'h0;
assign r_ram[921]= 7'h0;
assign r_ram[922]= 7'h0;
assign r_ram[923]= 7'h0;
assign r_ram[924]= 7'h11;
assign r_ram[925]= 7'h0;
assign r_ram[926]= 7'h0;
assign r_ram[927]= 7'h0;
assign r_ram[928]= 7'h0;
assign r_ram[929]= 7'h0;
assign r_ram[930]= 7'h0;
assign r_ram[931]= 7'h0;
assign r_ram[932]= 7'h0;
assign r_ram[933]= 7'h0;
assign r_ram[934]= 7'h0;
assign r_ram[935]= 7'h0;
assign r_ram[936]= 7'h0;
assign r_ram[937]= 7'h0;
assign r_ram[938]= 7'h0;
assign r_ram[939]= 7'h2;
assign r_ram[940]= 7'h0;
assign r_ram[941]= 7'h0;
assign r_ram[942]= 7'h0;
assign r_ram[943]= 7'h4;
assign r_ram[944]= 7'h8;
assign r_ram[945]= 7'h0;
assign r_ram[946]= 7'h0;
assign r_ram[947]= 7'h0;
assign r_ram[948]= 7'h0;
assign r_ram[949]= 7'h0;
assign r_ram[950]= 7'h0;
assign r_ram[951]= 7'h0;
assign r_ram[952]= 7'h0;
assign r_ram[953]= 7'h21;
assign r_ram[954]= 7'h0;
assign r_ram[955]= 7'h0;
assign r_ram[956]= 7'h0;
assign r_ram[957]= 7'h0;
assign r_ram[958]= 7'h0;
assign r_ram[959]= 7'h0;
assign r_ram[960]= 7'h0;
assign r_ram[961]= 7'h0;
assign r_ram[962]= 7'h0;
assign r_ram[963]= 7'h0;
assign r_ram[964]= 7'h0;
assign r_ram[965]= 7'h0;
assign r_ram[966]= 7'h0;
assign r_ram[967]= 7'h0;
assign r_ram[968]= 7'h0;
assign r_ram[969]= 7'h0;
assign r_ram[970]= 7'h0;
assign r_ram[971]= 7'h2;
assign r_ram[972]= 7'h0;
assign r_ram[973]= 7'h0;
assign r_ram[974]= 7'h0;
assign r_ram[975]= 7'h0;
assign r_ram[976]= 7'h0;
assign r_ram[977]= 7'h0;
assign r_ram[978]= 7'h0;
assign r_ram[979]= 7'h4;
assign r_ram[980]= 7'h0;
assign r_ram[981]= 7'h0;
assign r_ram[982]= 7'h0;
assign r_ram[983]= 7'h0;
assign r_ram[984]= 7'h8;
assign r_ram[985]= 7'h0;
assign r_ram[986]= 7'h41;
assign r_ram[987]= 7'h0;
assign r_ram[988]= 7'h0;
assign r_ram[989]= 7'h0;
assign r_ram[990]= 7'h0;
assign r_ram[991]= 7'h0;
assign r_ram[992]= 7'h0;
assign r_ram[993]= 7'h0;
assign r_ram[994]= 7'h0;
assign r_ram[995]= 7'h0;
assign r_ram[996]= 7'hc;
assign r_ram[997]= 7'h0;
assign r_ram[998]= 7'h0;
assign r_ram[999]= 7'h0;
assign r_ram[1000]= 7'h0;
assign r_ram[1001]= 7'h2;
assign r_ram[1002]= 7'h0;
assign r_ram[1003]= 7'h0;
assign r_ram[1004]= 7'h0;
assign r_ram[1005]= 7'h0;
assign r_ram[1006]= 7'h0;
assign r_ram[1007]= 7'h0;
assign r_ram[1008]= 7'h0;
assign r_ram[1009]= 7'h0;
assign r_ram[1010]= 7'h0;
assign r_ram[1011]= 7'h0;
assign r_ram[1012]= 7'h0;
assign r_ram[1013]= 7'h11;
assign r_ram[1014]= 7'h0;
assign r_ram[1015]= 7'h0;
assign r_ram[1016]= 7'h0;
assign r_ram[1017]= 7'h0;
assign r_ram[1018]= 7'h0;
assign r_ram[1019]= 7'h0;
assign r_ram[1020]= 7'h0;
assign r_ram[1021]= 7'h0;
assign r_ram[1022]= 7'h0;
assign r_ram[1023]= 7'h0;
assign r_ram[1024]= 7'h0;
assign r_ram[1025]= 7'h0;
assign r_ram[1026]= 7'h0;
assign r_ram[1027]= 7'h0;
assign r_ram[1028]= 7'h0;
assign r_ram[1029]= 7'h0;
assign r_ram[1030]= 7'h2;
assign r_ram[1031]= 7'h0;
assign r_ram[1032]= 7'h0;
assign r_ram[1033]= 7'h0;
assign r_ram[1034]= 7'h0;
assign r_ram[1035]= 7'h0;
assign r_ram[1036]= 7'h4;
assign r_ram[1037]= 7'h0;
assign r_ram[1038]= 7'h0;
assign r_ram[1039]= 7'h8;
assign r_ram[1040]= 7'h0;
assign r_ram[1041]= 7'h0;
assign r_ram[1042]= 7'h0;
assign r_ram[1043]= 7'h0;
assign r_ram[1044]= 7'h0;
assign r_ram[1045]= 7'h21;
assign r_ram[1046]= 7'h0;
assign r_ram[1047]= 7'h0;
assign r_ram[1048]= 7'h0;
assign r_ram[1049]= 7'h0;
assign r_ram[1050]= 7'h0;
assign r_ram[1051]= 7'h0;
assign r_ram[1052]= 7'h0;
assign r_ram[1053]= 7'h0;
assign r_ram[1054]= 7'h0;
assign r_ram[1055]= 7'h0;
assign r_ram[1056]= 7'h0;
assign r_ram[1057]= 7'h0;
assign r_ram[1058]= 7'h0;
assign r_ram[1059]= 7'h0;
assign r_ram[1060]= 7'h2;
assign r_ram[1061]= 7'h0;
assign r_ram[1062]= 7'h0;
assign r_ram[1063]= 7'h0;
assign r_ram[1064]= 7'h0;
assign r_ram[1065]= 7'h0;
assign r_ram[1066]= 7'h0;
assign r_ram[1067]= 7'h0;
assign r_ram[1068]= 7'h0;
assign r_ram[1069]= 7'h0;
assign r_ram[1070]= 7'h4;
assign r_ram[1071]= 7'h0;
assign r_ram[1072]= 7'h0;
assign r_ram[1073]= 7'h8;
assign r_ram[1074]= 7'h0;
assign r_ram[1075]= 7'h0;
assign r_ram[1076]= 7'h41;
assign r_ram[1077]= 7'h0;
assign r_ram[1078]= 7'h0;
assign r_ram[1079]= 7'h0;
assign r_ram[1080]= 7'h0;
assign r_ram[1081]= 7'h0;
assign r_ram[1082]= 7'h0;
assign r_ram[1083]= 7'h0;
assign r_ram[1084]= 7'h0;
assign r_ram[1085]= 7'hc;
assign r_ram[1086]= 7'h0;
assign r_ram[1087]= 7'h0;
assign r_ram[1088]= 7'h0;
assign r_ram[1089]= 7'h0;
assign r_ram[1090]= 7'h2;
assign r_ram[1091]= 7'h0;
assign r_ram[1092]= 7'h0;
assign r_ram[1093]= 7'h0;
assign r_ram[1094]= 7'h0;
assign r_ram[1095]= 7'h0;
assign r_ram[1096]= 7'h0;
assign r_ram[1097]= 7'h0;
assign r_ram[1098]= 7'h0;
assign r_ram[1099]= 7'h0;
assign r_ram[1100]= 7'h0;
assign r_ram[1101]= 7'h0;
assign r_ram[1102]= 7'h0;
assign r_ram[1103]= 7'h11;
assign r_ram[1104]= 7'h0;
assign r_ram[1105]= 7'h0;
assign r_ram[1106]= 7'h0;
assign r_ram[1107]= 7'h0;
assign r_ram[1108]= 7'h0;
assign r_ram[1109]= 7'h0;
assign r_ram[1110]= 7'h0;
assign r_ram[1111]= 7'h0;
assign r_ram[1112]= 7'h0;
assign r_ram[1113]= 7'h0;
assign r_ram[1114]= 7'h0;
assign r_ram[1115]= 7'h0;
assign r_ram[1116]= 7'h0;
assign r_ram[1117]= 7'h0;
assign r_ram[1118]= 7'h0;
assign r_ram[1119]= 7'h2;
assign r_ram[1120]= 7'h0;
assign r_ram[1121]= 7'h0;
assign r_ram[1122]= 7'h0;
assign r_ram[1123]= 7'h0;
assign r_ram[1124]= 7'h8;
assign r_ram[1125]= 7'h4;
assign r_ram[1126]= 7'h0;
assign r_ram[1127]= 7'h0;
assign r_ram[1128]= 7'h0;
assign r_ram[1129]= 7'h0;
assign r_ram[1130]= 7'h0;
assign r_ram[1131]= 7'h0;
assign r_ram[1132]= 7'h0;
assign r_ram[1133]= 7'h0;
assign r_ram[1134]= 7'h0;
assign r_ram[1135]= 7'h21;
assign r_ram[1136]= 7'h0;
assign r_ram[1137]= 7'h0;
assign r_ram[1138]= 7'h0;
assign r_ram[1139]= 7'h0;
assign r_ram[1140]= 7'h0;
assign r_ram[1141]= 7'h0;
assign r_ram[1142]= 7'h0;
assign r_ram[1143]= 7'h0;
assign r_ram[1144]= 7'h0;
assign r_ram[1145]= 7'h0;
assign r_ram[1146]= 7'h0;
assign r_ram[1147]= 7'h0;
assign r_ram[1148]= 7'h0;
assign r_ram[1149]= 7'h0;
assign r_ram[1150]= 7'h2;
assign r_ram[1151]= 7'h0;
assign r_ram[1152]= 7'h0;
assign r_ram[1153]= 7'h0;
assign r_ram[1154]= 7'h0;
assign r_ram[1155]= 7'h0;
assign r_ram[1156]= 7'h0;
assign r_ram[1157]= 7'h0;
assign r_ram[1158]= 7'h0;
assign r_ram[1159]= 7'h0;
assign r_ram[1160]= 7'h0;
assign r_ram[1161]= 7'h4;
assign r_ram[1162]= 7'h0;
assign r_ram[1163]= 7'h0;
assign r_ram[1164]= 7'h0;
assign r_ram[1165]= 7'h8;
assign r_ram[1166]= 7'h0;
assign r_ram[1167]= 7'h41;
assign r_ram[1168]= 7'h0;
assign r_ram[1169]= 7'h0;
assign r_ram[1170]= 7'h0;
assign r_ram[1171]= 7'h0;
assign r_ram[1172]= 7'h0;
assign r_ram[1173]= 7'h0;
assign r_ram[1174]= 7'h4;
assign r_ram[1175]= 7'h8;
assign r_ram[1176]= 7'h0;
assign r_ram[1177]= 7'h0;
assign r_ram[1178]= 7'h0;
assign r_ram[1179]= 7'h0;
assign r_ram[1180]= 7'h2;
assign r_ram[1181]= 7'h0;
assign r_ram[1182]= 7'h0;
assign r_ram[1183]= 7'h0;
assign r_ram[1184]= 7'h0;
assign r_ram[1185]= 7'h0;
assign r_ram[1186]= 7'h0;
assign r_ram[1187]= 7'h0;
assign r_ram[1188]= 7'h0;
assign r_ram[1189]= 7'h0;
assign r_ram[1190]= 7'h0;
assign r_ram[1191]= 7'h0;
assign r_ram[1192]= 7'h11;
assign r_ram[1193]= 7'h0;
assign r_ram[1194]= 7'h0;
assign r_ram[1195]= 7'h0;
assign r_ram[1196]= 7'h0;
assign r_ram[1197]= 7'h0;
assign r_ram[1198]= 7'h0;
assign r_ram[1199]= 7'h0;
assign r_ram[1200]= 7'h0;
assign r_ram[1201]= 7'h0;
assign r_ram[1202]= 7'h0;
assign r_ram[1203]= 7'h0;
assign r_ram[1204]= 7'h0;
assign r_ram[1205]= 7'h0;
assign r_ram[1206]= 7'h0;
assign r_ram[1207]= 7'h0;
assign r_ram[1208]= 7'h0;
assign r_ram[1209]= 7'h0;
assign r_ram[1210]= 7'h2;
assign r_ram[1211]= 7'h0;
assign r_ram[1212]= 7'h0;
assign r_ram[1213]= 7'h0;
assign r_ram[1214]= 7'h0;
assign r_ram[1215]= 7'h0;
assign r_ram[1216]= 7'h0;
assign r_ram[1217]= 7'h0;
assign r_ram[1218]= 7'hc;
assign r_ram[1219]= 7'h0;
assign r_ram[1220]= 7'h0;
assign r_ram[1221]= 7'h0;
assign r_ram[1222]= 7'h0;
assign r_ram[1223]= 7'h0;
assign r_ram[1224]= 7'h0;
assign r_ram[1225]= 7'h21;
assign r_ram[1226]= 7'h0;
assign r_ram[1227]= 7'h0;
assign r_ram[1228]= 7'h0;
assign r_ram[1229]= 7'h0;
assign r_ram[1230]= 7'h0;
assign r_ram[1231]= 7'h0;
assign r_ram[1232]= 7'h0;
assign r_ram[1233]= 7'h0;
assign r_ram[1234]= 7'h0;
assign r_ram[1235]= 7'h0;
assign r_ram[1236]= 7'h0;
assign r_ram[1237]= 7'h0;
assign r_ram[1238]= 7'h0;
assign r_ram[1239]= 7'h0;
assign r_ram[1240]= 7'h2;
assign r_ram[1241]= 7'h0;
assign r_ram[1242]= 7'h0;
assign r_ram[1243]= 7'h0;
assign r_ram[1244]= 7'h0;
assign r_ram[1245]= 7'h0;
assign r_ram[1246]= 7'h0;
assign r_ram[1247]= 7'h0;
assign r_ram[1248]= 7'h0;
assign r_ram[1249]= 7'h4;
assign r_ram[1250]= 7'h0;
assign r_ram[1251]= 7'h0;
assign r_ram[1252]= 7'h0;
assign r_ram[1253]= 7'h0;
assign r_ram[1254]= 7'h8;
assign r_ram[1255]= 7'h41;
assign r_ram[1256]= 7'h0;
assign r_ram[1257]= 7'h0;
assign r_ram[1258]= 7'h0;
assign r_ram[1259]= 7'h0;
assign r_ram[1260]= 7'h0;
assign r_ram[1261]= 7'h0;
assign r_ram[1262]= 7'h0;
assign r_ram[1263]= 7'h0;
assign r_ram[1264]= 7'h4;
assign r_ram[1265]= 7'h0;
assign r_ram[1266]= 7'h8;
assign r_ram[1267]= 7'h0;
assign r_ram[1268]= 7'h0;
assign r_ram[1269]= 7'h0;
assign r_ram[1270]= 7'h0;
assign r_ram[1271]= 7'h0;
assign r_ram[1272]= 7'h2;
assign r_ram[1273]= 7'h0;
assign r_ram[1274]= 7'h0;
assign r_ram[1275]= 7'h0;
assign r_ram[1276]= 7'h0;
assign r_ram[1277]= 7'h0;
assign r_ram[1278]= 7'h0;
assign r_ram[1279]= 7'h0;
assign r_ram[1280]= 7'h0;
assign r_ram[1281]= 7'h0;
assign r_ram[1282]= 7'h0;
assign r_ram[1283]= 7'h0;
assign r_ram[1284]= 7'h0;
assign r_ram[1285]= 7'h11;
assign r_ram[1286]= 7'h0;
assign r_ram[1287]= 7'h0;
assign r_ram[1288]= 7'h0;
assign r_ram[1289]= 7'h0;
assign r_ram[1290]= 7'h0;
assign r_ram[1291]= 7'h0;
assign r_ram[1292]= 7'h0;
assign r_ram[1293]= 7'h0;
assign r_ram[1294]= 7'h0;
assign r_ram[1295]= 7'h0;
assign r_ram[1296]= 7'h0;
assign r_ram[1297]= 7'h0;
assign r_ram[1298]= 7'h0;
assign r_ram[1299]= 7'h0;
assign r_ram[1300]= 7'h2;
assign r_ram[1301]= 7'h0;
assign r_ram[1302]= 7'h0;
assign r_ram[1303]= 7'h0;
assign r_ram[1304]= 7'h4;
assign r_ram[1305]= 7'h0;
assign r_ram[1306]= 7'h0;
assign r_ram[1307]= 7'h8;
assign r_ram[1308]= 7'h0;
assign r_ram[1309]= 7'h0;
assign r_ram[1310]= 7'h0;
assign r_ram[1311]= 7'h0;
assign r_ram[1312]= 7'h0;
assign r_ram[1313]= 7'h0;
assign r_ram[1314]= 7'h21;
assign r_ram[1315]= 7'h0;
assign r_ram[1316]= 7'h0;
assign r_ram[1317]= 7'h0;
assign r_ram[1318]= 7'h0;
assign r_ram[1319]= 7'h0;
assign r_ram[1320]= 7'h0;
assign r_ram[1321]= 7'h0;
assign r_ram[1322]= 7'h0;
assign r_ram[1323]= 7'h0;
assign r_ram[1324]= 7'h0;
assign r_ram[1325]= 7'h0;
assign r_ram[1326]= 7'h0;
assign r_ram[1327]= 7'h0;
assign r_ram[1328]= 7'h0;
assign r_ram[1329]= 7'h0;
assign r_ram[1330]= 7'h2;
assign r_ram[1331]= 7'h0;
assign r_ram[1332]= 7'h0;
assign r_ram[1333]= 7'h0;
assign r_ram[1334]= 7'h0;
assign r_ram[1335]= 7'h0;
assign r_ram[1336]= 7'h0;
assign r_ram[1337]= 7'h0;
assign r_ram[1338]= 7'h0;
assign r_ram[1339]= 7'h4;
assign r_ram[1340]= 7'h0;
assign r_ram[1341]= 7'h0;
assign r_ram[1342]= 7'h0;
assign r_ram[1343]= 7'h0;
assign r_ram[1344]= 7'h0;
assign r_ram[1345]= 7'h1;
assign r_ram[1346]= 7'h0;
assign r_ram[1347]= 7'h0;
assign r_ram[1348]= 7'h48;
assign r_ram[1349]= 7'h0;
assign r_ram[1350]= 7'h0;
assign r_ram[1351]= 7'h0;
assign r_ram[1352]= 7'h0;
assign r_ram[1353]= 7'h0;
assign r_ram[1354]= 7'h0;
assign r_ram[1355]= 7'h0;
assign r_ram[1356]= 7'h4;
assign r_ram[1357]= 7'h0;
assign r_ram[1358]= 7'h8;
assign r_ram[1359]= 7'h0;
assign r_ram[1360]= 7'h0;
assign r_ram[1361]= 7'h0;
assign r_ram[1362]= 7'h2;
assign r_ram[1363]= 7'h0;
assign r_ram[1364]= 7'h0;
assign r_ram[1365]= 7'h0;
assign r_ram[1366]= 7'h0;
assign r_ram[1367]= 7'h0;
assign r_ram[1368]= 7'h0;
assign r_ram[1369]= 7'h0;
assign r_ram[1370]= 7'h0;
assign r_ram[1371]= 7'h0;
assign r_ram[1372]= 7'h0;
assign r_ram[1373]= 7'h0;
assign r_ram[1374]= 7'h0;
assign r_ram[1375]= 7'h11;
assign r_ram[1376]= 7'h0;
assign r_ram[1377]= 7'h0;
assign r_ram[1378]= 7'h0;
assign r_ram[1379]= 7'h0;
assign r_ram[1380]= 7'h0;
assign r_ram[1381]= 7'h0;
assign r_ram[1382]= 7'h0;
assign r_ram[1383]= 7'h0;
assign r_ram[1384]= 7'h0;
assign r_ram[1385]= 7'h0;
assign r_ram[1386]= 7'h0;
assign r_ram[1387]= 7'h0;
assign r_ram[1388]= 7'h0;
assign r_ram[1389]= 7'h0;
assign r_ram[1390]= 7'h2;
assign r_ram[1391]= 7'h0;
assign r_ram[1392]= 7'h0;
assign r_ram[1393]= 7'h0;
assign r_ram[1394]= 7'h0;
assign r_ram[1395]= 7'h0;
assign r_ram[1396]= 7'h0;
assign r_ram[1397]= 7'h4;
assign r_ram[1398]= 7'h8;
assign r_ram[1399]= 7'h0;
assign r_ram[1400]= 7'h0;
assign r_ram[1401]= 7'h0;
assign r_ram[1402]= 7'h0;
assign r_ram[1403]= 7'h0;
assign r_ram[1404]= 7'h0;
assign r_ram[1405]= 7'h0;
assign r_ram[1406]= 7'h21;
assign r_ram[1407]= 7'h0;
assign r_ram[1408]= 7'h0;
assign r_ram[1409]= 7'h0;
assign r_ram[1410]= 7'h0;
assign r_ram[1411]= 7'h0;
assign r_ram[1412]= 7'h0;
assign r_ram[1413]= 7'h0;
assign r_ram[1414]= 7'h0;
assign r_ram[1415]= 7'h0;
assign r_ram[1416]= 7'h0;
assign r_ram[1417]= 7'h0;
assign r_ram[1418]= 7'h0;
assign r_ram[1419]= 7'h0;
assign r_ram[1420]= 7'h0;
assign r_ram[1421]= 7'h2;
assign r_ram[1422]= 7'h0;
assign r_ram[1423]= 7'h0;
assign r_ram[1424]= 7'h0;
assign r_ram[1425]= 7'h0;
assign r_ram[1426]= 7'h0;
assign r_ram[1427]= 7'h0;
assign r_ram[1428]= 7'h0;
assign r_ram[1429]= 7'h0;
assign r_ram[1430]= 7'h4;
assign r_ram[1431]= 7'h0;
assign r_ram[1432]= 7'h0;
assign r_ram[1433]= 7'h0;
assign r_ram[1434]= 7'h0;
assign r_ram[1435]= 7'h0;
assign r_ram[1436]= 7'h1;
assign r_ram[1437]= 7'h48;
assign r_ram[1438]= 7'h0;
assign r_ram[1439]= 7'h0;
assign r_ram[1440]= 7'h0;
assign r_ram[1441]= 7'h0;
assign r_ram[1442]= 7'h0;
assign r_ram[1443]= 7'h0;
assign r_ram[1444]= 7'h0;
assign r_ram[1445]= 7'h4;
assign r_ram[1446]= 7'h0;
assign r_ram[1447]= 7'h0;
assign r_ram[1448]= 7'h8;
assign r_ram[1449]= 7'h0;
assign r_ram[1450]= 7'h0;
assign r_ram[1451]= 7'h2;
assign r_ram[1452]= 7'h0;
assign r_ram[1453]= 7'h0;
assign r_ram[1454]= 7'h0;
assign r_ram[1455]= 7'h0;
assign r_ram[1456]= 7'h0;
assign r_ram[1457]= 7'h0;
assign r_ram[1458]= 7'h0;
assign r_ram[1459]= 7'h0;
assign r_ram[1460]= 7'h0;
assign r_ram[1461]= 7'h0;
assign r_ram[1462]= 7'h0;
assign r_ram[1463]= 7'h0;
assign r_ram[1464]= 7'h11;
assign r_ram[1465]= 7'h0;
assign r_ram[1466]= 7'h0;
assign r_ram[1467]= 7'h0;
assign r_ram[1468]= 7'h0;
assign r_ram[1469]= 7'h0;
assign r_ram[1470]= 7'h0;
assign r_ram[1471]= 7'h0;
assign r_ram[1472]= 7'h0;
assign r_ram[1473]= 7'h0;
assign r_ram[1474]= 7'h0;
assign r_ram[1475]= 7'h0;
assign r_ram[1476]= 7'h0;
assign r_ram[1477]= 7'h0;
assign r_ram[1478]= 7'h0;
assign r_ram[1479]= 7'h0;
assign r_ram[1480]= 7'h2;
assign r_ram[1481]= 7'h0;
assign r_ram[1482]= 7'h0;
assign r_ram[1483]= 7'h0;
assign r_ram[1484]= 7'h0;
assign r_ram[1485]= 7'h0;
assign r_ram[1486]= 7'h0;
assign r_ram[1487]= 7'h4;
assign r_ram[1488]= 7'h0;
assign r_ram[1489]= 7'h8;
assign r_ram[1490]= 7'h0;
assign r_ram[1491]= 7'h0;
assign r_ram[1492]= 7'h0;
assign r_ram[1493]= 7'h0;
assign r_ram[1494]= 7'h21;
assign r_ram[1495]= 7'h0;
assign r_ram[1496]= 7'h0;
assign r_ram[1497]= 7'h0;
assign r_ram[1498]= 7'h0;
assign r_ram[1499]= 7'h0;
assign r_ram[1500]= 7'h0;
assign r_ram[1501]= 7'h0;
assign r_ram[1502]= 7'h0;
assign r_ram[1503]= 7'h0;
assign r_ram[1504]= 7'h0;
assign r_ram[1505]= 7'h0;
assign r_ram[1506]= 7'h0;
assign r_ram[1507]= 7'h0;
assign r_ram[1508]= 7'h0;
assign r_ram[1509]= 7'h0;
assign r_ram[1510]= 7'h2;
assign r_ram[1511]= 7'h0;
assign r_ram[1512]= 7'h0;
assign r_ram[1513]= 7'h0;
assign r_ram[1514]= 7'h0;
assign r_ram[1515]= 7'h0;
assign r_ram[1516]= 7'h0;
assign r_ram[1517]= 7'h0;
assign r_ram[1518]= 7'h0;
assign r_ram[1519]= 7'h0;
assign r_ram[1520]= 7'h0;
assign r_ram[1521]= 7'h4;
assign r_ram[1522]= 7'h8;
assign r_ram[1523]= 7'h0;
assign r_ram[1524]= 7'h0;
assign r_ram[1525]= 7'h0;
assign r_ram[1526]= 7'h41;
assign r_ram[1527]= 7'h0;
assign r_ram[1528]= 7'h0;
assign r_ram[1529]= 7'h0;
assign r_ram[1530]= 7'h0;
assign r_ram[1531]= 7'h0;
assign r_ram[1532]= 7'h0;
assign r_ram[1533]= 7'h0;
assign r_ram[1534]= 7'h0;
assign r_ram[1535]= 7'h4;
assign r_ram[1536]= 7'h0;
assign r_ram[1537]= 7'h8;
assign r_ram[1538]= 7'h0;
assign r_ram[1539]= 7'h0;
assign r_ram[1540]= 7'h0;
assign r_ram[1541]= 7'h2;
assign r_ram[1542]= 7'h0;
assign r_ram[1543]= 7'h0;
assign r_ram[1544]= 7'h0;
assign r_ram[1545]= 7'h0;
assign r_ram[1546]= 7'h0;
assign r_ram[1547]= 7'h0;
assign r_ram[1548]= 7'h0;
assign r_ram[1549]= 7'h0;
assign r_ram[1550]= 7'h0;
assign r_ram[1551]= 7'h0;
assign r_ram[1552]= 7'h0;
assign r_ram[1553]= 7'h11;
assign r_ram[1554]= 7'h0;
assign r_ram[1555]= 7'h0;
assign r_ram[1556]= 7'h0;
assign r_ram[1557]= 7'h0;
assign r_ram[1558]= 7'h0;
assign r_ram[1559]= 7'h0;
assign r_ram[1560]= 7'h0;
assign r_ram[1561]= 7'h0;
assign r_ram[1562]= 7'h0;
assign r_ram[1563]= 7'h0;
assign r_ram[1564]= 7'h0;
assign r_ram[1565]= 7'h0;
assign r_ram[1566]= 7'h0;
assign r_ram[1567]= 7'h0;
assign r_ram[1568]= 7'h0;
assign r_ram[1569]= 7'h0;
assign r_ram[1570]= 7'h2;
assign r_ram[1571]= 7'h0;
assign r_ram[1572]= 7'h0;
assign r_ram[1573]= 7'h0;
assign r_ram[1574]= 7'h8;
assign r_ram[1575]= 7'h4;
assign r_ram[1576]= 7'h0;
assign r_ram[1577]= 7'h0;
assign r_ram[1578]= 7'h0;
assign r_ram[1579]= 7'h0;
assign r_ram[1580]= 7'h0;
assign r_ram[1581]= 7'h0;
assign r_ram[1582]= 7'h0;
assign r_ram[1583]= 7'h0;
assign r_ram[1584]= 7'h0;
assign r_ram[1585]= 7'h21;
assign r_ram[1586]= 7'h0;
assign r_ram[1587]= 7'h0;
assign r_ram[1588]= 7'h0;
assign r_ram[1589]= 7'h0;
assign r_ram[1590]= 7'h0;
assign r_ram[1591]= 7'h0;
assign r_ram[1592]= 7'h0;
assign r_ram[1593]= 7'h0;
assign r_ram[1594]= 7'h0;
assign r_ram[1595]= 7'h0;
assign r_ram[1596]= 7'h0;
assign r_ram[1597]= 7'h0;
assign r_ram[1598]= 7'h0;
assign r_ram[1599]= 7'h0;
assign r_ram[1600]= 7'h0;
assign r_ram[1601]= 7'h2;
assign r_ram[1602]= 7'h0;
assign r_ram[1603]= 7'h0;
assign r_ram[1604]= 7'h0;
assign r_ram[1605]= 7'h0;
assign r_ram[1606]= 7'h0;
assign r_ram[1607]= 7'h0;
assign r_ram[1608]= 7'h0;
assign r_ram[1609]= 7'h0;
assign r_ram[1610]= 7'h0;
assign r_ram[1611]= 7'h0;
assign r_ram[1612]= 7'h0;
assign r_ram[1613]= 7'h0;
assign r_ram[1614]= 7'h0;
assign r_ram[1615]= 7'h4;
assign r_ram[1616]= 7'h8;
assign r_ram[1617]= 7'h0;
assign r_ram[1618]= 7'h41;
assign r_ram[1619]= 7'h0;
assign r_ram[1620]= 7'h0;
assign r_ram[1621]= 7'h0;
assign r_ram[1622]= 7'h0;
assign r_ram[1623]= 7'h0;
assign r_ram[1624]= 7'h0;
assign r_ram[1625]= 7'h0;
assign r_ram[1626]= 7'h4;
assign r_ram[1627]= 7'h8;
assign r_ram[1628]= 7'h0;
assign r_ram[1629]= 7'h0;
assign r_ram[1630]= 7'h0;
assign r_ram[1631]= 7'h2;
assign r_ram[1632]= 7'h0;
assign r_ram[1633]= 7'h0;
assign r_ram[1634]= 7'h0;
assign r_ram[1635]= 7'h0;
assign r_ram[1636]= 7'h0;
assign r_ram[1637]= 7'h0;
assign r_ram[1638]= 7'h0;
assign r_ram[1639]= 7'h0;
assign r_ram[1640]= 7'h0;
assign r_ram[1641]= 7'h0;
assign r_ram[1642]= 7'h0;
assign r_ram[1643]= 7'h0;
assign r_ram[1644]= 7'h0;
assign r_ram[1645]= 7'h11;
assign r_ram[1646]= 7'h0;
assign r_ram[1647]= 7'h0;
assign r_ram[1648]= 7'h0;
assign r_ram[1649]= 7'h0;
assign r_ram[1650]= 7'h0;
assign r_ram[1651]= 7'h0;
assign r_ram[1652]= 7'h0;
assign r_ram[1653]= 7'h0;
assign r_ram[1654]= 7'h0;
assign r_ram[1655]= 7'h0;
assign r_ram[1656]= 7'h0;
assign r_ram[1657]= 7'h0;
assign r_ram[1658]= 7'h0;
assign r_ram[1659]= 7'h2;
assign r_ram[1660]= 7'h0;
assign r_ram[1661]= 7'h0;
assign r_ram[1662]= 7'h0;
assign r_ram[1663]= 7'h0;
assign r_ram[1664]= 7'h0;
assign r_ram[1665]= 7'h0;
assign r_ram[1666]= 7'h0;
assign r_ram[1667]= 7'h4;
assign r_ram[1668]= 7'h0;
assign r_ram[1669]= 7'h8;
assign r_ram[1670]= 7'h0;
assign r_ram[1671]= 7'h0;
assign r_ram[1672]= 7'h0;
assign r_ram[1673]= 7'h0;
assign r_ram[1674]= 7'h0;
assign r_ram[1675]= 7'h0;
assign r_ram[1676]= 7'h21;
assign r_ram[1677]= 7'h0;
assign r_ram[1678]= 7'h0;
assign r_ram[1679]= 7'h0;
assign r_ram[1680]= 7'h0;
assign r_ram[1681]= 7'h0;
assign r_ram[1682]= 7'h0;
assign r_ram[1683]= 7'h0;
assign r_ram[1684]= 7'h0;
assign r_ram[1685]= 7'h0;
assign r_ram[1686]= 7'h0;
assign r_ram[1687]= 7'h0;
assign r_ram[1688]= 7'h0;
assign r_ram[1689]= 7'h0;
assign r_ram[1690]= 7'h2;
assign r_ram[1691]= 7'h0;
assign r_ram[1692]= 7'h0;
assign r_ram[1693]= 7'h0;
assign r_ram[1694]= 7'h0;
assign r_ram[1695]= 7'h0;
assign r_ram[1696]= 7'h0;
assign r_ram[1697]= 7'h0;
assign r_ram[1698]= 7'h0;
assign r_ram[1699]= 7'h0;
assign r_ram[1700]= 7'h0;
assign r_ram[1701]= 7'h0;
assign r_ram[1702]= 7'h0;
assign r_ram[1703]= 7'h0;
assign r_ram[1704]= 7'h0;
assign r_ram[1705]= 7'h0;
assign r_ram[1706]= 7'h4;
assign r_ram[1707]= 7'h8;
assign r_ram[1708]= 7'h41;
assign r_ram[1709]= 7'h0;
assign r_ram[1710]= 7'h0;
assign r_ram[1711]= 7'h0;
assign r_ram[1712]= 7'h0;
assign r_ram[1713]= 7'h0;
assign r_ram[1714]= 7'h0;
assign r_ram[1715]= 7'h0;
assign r_ram[1716]= 7'h4;
assign r_ram[1717]= 7'h8;
assign r_ram[1718]= 7'h0;
assign r_ram[1719]= 7'h0;
assign r_ram[1720]= 7'h0;
assign r_ram[1721]= 7'h2;
assign r_ram[1722]= 7'h0;
assign r_ram[1723]= 7'h0;
assign r_ram[1724]= 7'h0;
assign r_ram[1725]= 7'h0;
assign r_ram[1726]= 7'h0;
assign r_ram[1727]= 7'h0;
assign r_ram[1728]= 7'h0;
assign r_ram[1729]= 7'h0;
assign r_ram[1730]= 7'h0;
assign r_ram[1731]= 7'h0;
assign r_ram[1732]= 7'h0;
assign r_ram[1733]= 7'h11;
assign r_ram[1734]= 7'h0;
assign r_ram[1735]= 7'h0;
assign r_ram[1736]= 7'h0;
assign r_ram[1737]= 7'h0;
assign r_ram[1738]= 7'h0;
assign r_ram[1739]= 7'h0;
assign r_ram[1740]= 7'h0;
assign r_ram[1741]= 7'h0;
assign r_ram[1742]= 7'h0;
assign r_ram[1743]= 7'h0;
assign r_ram[1744]= 7'h0;
assign r_ram[1745]= 7'h0;
assign r_ram[1746]= 7'h0;
assign r_ram[1747]= 7'h0;
assign r_ram[1748]= 7'h0;
assign r_ram[1749]= 7'h0;
assign r_ram[1750]= 7'h2;
assign r_ram[1751]= 7'h0;
assign r_ram[1752]= 7'h0;
assign r_ram[1753]= 7'h0;
assign r_ram[1754]= 7'h0;
assign r_ram[1755]= 7'hc;
assign r_ram[1756]= 7'h0;
assign r_ram[1757]= 7'h0;
assign r_ram[1758]= 7'h0;
assign r_ram[1759]= 7'h0;
assign r_ram[1760]= 7'h0;
assign r_ram[1761]= 7'h0;
assign r_ram[1762]= 7'h0;
assign r_ram[1763]= 7'h0;
assign r_ram[1764]= 7'h21;
assign r_ram[1765]= 7'h0;
assign r_ram[1766]= 7'h0;
assign r_ram[1767]= 7'h0;
assign r_ram[1768]= 7'h0;
assign r_ram[1769]= 7'h0;
assign r_ram[1770]= 7'h0;
assign r_ram[1771]= 7'h0;
assign r_ram[1772]= 7'h0;
assign r_ram[1773]= 7'h0;
assign r_ram[1774]= 7'h0;
assign r_ram[1775]= 7'h0;
assign r_ram[1776]= 7'h0;
assign r_ram[1777]= 7'h0;
assign r_ram[1778]= 7'h0;
assign r_ram[1779]= 7'h2;
assign r_ram[1780]= 7'h0;
assign r_ram[1781]= 7'h0;
assign r_ram[1782]= 7'h0;
assign r_ram[1783]= 7'h0;
assign r_ram[1784]= 7'h0;
assign r_ram[1785]= 7'h0;
assign r_ram[1786]= 7'h0;
assign r_ram[1787]= 7'h0;
assign r_ram[1788]= 7'h0;
assign r_ram[1789]= 7'hc;
assign r_ram[1790]= 7'h0;
assign r_ram[1791]= 7'h0;
assign r_ram[1792]= 7'h0;
assign r_ram[1793]= 7'h0;
assign r_ram[1794]= 7'h0;
assign r_ram[1795]= 7'h41;
assign r_ram[1796]= 7'h0;
assign r_ram[1797]= 7'h0;
assign r_ram[1798]= 7'h0;
assign r_ram[1799]= 7'h0;
assign r_ram[1800]= 7'h0;
assign r_ram[1801]= 7'h0;
assign r_ram[1802]= 7'h0;
assign r_ram[1803]= 7'h0;
assign r_ram[1804]= 7'h0;
assign r_ram[1805]= 7'h0;
assign r_ram[1806]= 7'hc;
assign r_ram[1807]= 7'h0;
assign r_ram[1808]= 7'h0;
assign r_ram[1809]= 7'h0;
assign r_ram[1810]= 7'h0;
assign r_ram[1811]= 7'h2;
assign r_ram[1812]= 7'h0;
assign r_ram[1813]= 7'h0;
assign r_ram[1814]= 7'h0;
assign r_ram[1815]= 7'h0;
assign r_ram[1816]= 7'h0;
assign r_ram[1817]= 7'h0;
assign r_ram[1818]= 7'h0;
assign r_ram[1819]= 7'h0;
assign r_ram[1820]= 7'h0;
assign r_ram[1821]= 7'h0;
assign r_ram[1822]= 7'h0;
assign r_ram[1823]= 7'h0;
assign r_ram[1824]= 7'h11;
assign r_ram[1825]= 7'h0;
assign r_ram[1826]= 7'h0;
assign r_ram[1827]= 7'h0;
assign r_ram[1828]= 7'h0;
assign r_ram[1829]= 7'h0;
assign r_ram[1830]= 7'h0;
assign r_ram[1831]= 7'h0;
assign r_ram[1832]= 7'h0;
assign r_ram[1833]= 7'h0;
assign r_ram[1834]= 7'h0;
assign r_ram[1835]= 7'h0;
assign r_ram[1836]= 7'h0;
assign r_ram[1837]= 7'h0;
assign r_ram[1838]= 7'h0;
assign r_ram[1839]= 7'h0;
assign r_ram[1840]= 7'h0;
assign r_ram[1841]= 7'h2;
assign r_ram[1842]= 7'h0;
assign r_ram[1843]= 7'h0;
assign r_ram[1844]= 7'h0;
assign r_ram[1845]= 7'h0;
assign r_ram[1846]= 7'h0;
assign r_ram[1847]= 7'h0;
assign r_ram[1848]= 7'h4;
assign r_ram[1849]= 7'h0;
assign r_ram[1850]= 7'h0;
assign r_ram[1851]= 7'h0;
assign r_ram[1852]= 7'h8;
assign r_ram[1853]= 7'h0;
assign r_ram[1854]= 7'h0;
assign r_ram[1855]= 7'h21;
assign r_ram[1856]= 7'h0;
assign r_ram[1857]= 7'h0;
assign r_ram[1858]= 7'h0;
assign r_ram[1859]= 7'h0;
assign r_ram[1860]= 7'h0;
assign r_ram[1861]= 7'h0;
assign r_ram[1862]= 7'h0;
assign r_ram[1863]= 7'h0;
assign r_ram[1864]= 7'h0;
assign r_ram[1865]= 7'h0;
assign r_ram[1866]= 7'h0;
assign r_ram[1867]= 7'h0;
assign r_ram[1868]= 7'h0;
assign r_ram[1869]= 7'h0;
assign r_ram[1870]= 7'h0;
assign r_ram[1871]= 7'h2;
assign r_ram[1872]= 7'h0;
assign r_ram[1873]= 7'h0;
assign r_ram[1874]= 7'h0;
assign r_ram[1875]= 7'h0;
assign r_ram[1876]= 7'h0;
assign r_ram[1877]= 7'h0;
assign r_ram[1878]= 7'h0;
assign r_ram[1879]= 7'h0;
assign r_ram[1880]= 7'h0;
assign r_ram[1881]= 7'h0;
assign r_ram[1882]= 7'h4;
assign r_ram[1883]= 7'h0;
assign r_ram[1884]= 7'h0;
assign r_ram[1885]= 7'h0;
assign r_ram[1886]= 7'h0;
assign r_ram[1887]= 7'h49;
assign r_ram[1888]= 7'h0;
assign r_ram[1889]= 7'h0;
assign r_ram[1890]= 7'h0;
assign r_ram[1891]= 7'h0;
assign r_ram[1892]= 7'h0;
assign r_ram[1893]= 7'h0;
assign r_ram[1894]= 7'h0;
assign r_ram[1895]= 7'h0;
assign r_ram[1896]= 7'h4;
assign r_ram[1897]= 7'h0;
assign r_ram[1898]= 7'h8;
assign r_ram[1899]= 7'h0;
assign r_ram[1900]= 7'h0;
assign r_ram[1901]= 7'h2;
assign r_ram[1902]= 7'h0;
assign r_ram[1903]= 7'h0;
assign r_ram[1904]= 7'h0;
assign r_ram[1905]= 7'h0;
assign r_ram[1906]= 7'h0;
assign r_ram[1907]= 7'h0;
assign r_ram[1908]= 7'h0;
assign r_ram[1909]= 7'h0;
assign r_ram[1910]= 7'h0;
assign r_ram[1911]= 7'h0;
assign r_ram[1912]= 7'h0;
assign r_ram[1913]= 7'h11;
assign r_ram[1914]= 7'h0;
assign r_ram[1915]= 7'h0;
assign r_ram[1916]= 7'h0;
assign r_ram[1917]= 7'h0;
assign r_ram[1918]= 7'h0;
assign r_ram[1919]= 7'h0;
assign r_ram[1920]= 7'h0;
assign r_ram[1921]= 7'h0;
assign r_ram[1922]= 7'h0;
assign r_ram[1923]= 7'h0;
assign r_ram[1924]= 7'h0;
assign r_ram[1925]= 7'h0;
assign r_ram[1926]= 7'h0;
assign r_ram[1927]= 7'h0;
assign r_ram[1928]= 7'h0;
assign r_ram[1929]= 7'h0;
assign r_ram[1930]= 7'h2;
assign r_ram[1931]= 7'h0;
assign r_ram[1932]= 7'h0;
assign r_ram[1933]= 7'h0;
assign r_ram[1934]= 7'h0;
assign r_ram[1935]= 7'h4;
assign r_ram[1936]= 7'h0;
assign r_ram[1937]= 7'h8;
assign r_ram[1938]= 7'h0;
assign r_ram[1939]= 7'h0;
assign r_ram[1940]= 7'h0;
assign r_ram[1941]= 7'h0;
assign r_ram[1942]= 7'h0;
assign r_ram[1943]= 7'h0;
assign r_ram[1944]= 7'h0;
assign r_ram[1945]= 7'h21;
assign r_ram[1946]= 7'h0;
assign r_ram[1947]= 7'h0;
assign r_ram[1948]= 7'h0;
assign r_ram[1949]= 7'h0;
assign r_ram[1950]= 7'h0;
assign r_ram[1951]= 7'h0;
assign r_ram[1952]= 7'h0;
assign r_ram[1953]= 7'h0;
assign r_ram[1954]= 7'h0;
assign r_ram[1955]= 7'h0;
assign r_ram[1956]= 7'h0;
assign r_ram[1957]= 7'h0;
assign r_ram[1958]= 7'h0;
assign r_ram[1959]= 7'h0;
assign r_ram[1960]= 7'h2;
assign r_ram[1961]= 7'h0;
assign r_ram[1962]= 7'h0;
assign r_ram[1963]= 7'h0;
assign r_ram[1964]= 7'h0;
assign r_ram[1965]= 7'h0;
assign r_ram[1966]= 7'h0;
assign r_ram[1967]= 7'h0;
assign r_ram[1968]= 7'h0;
assign r_ram[1969]= 7'h4;
assign r_ram[1970]= 7'h0;
assign r_ram[1971]= 7'h0;
assign r_ram[1972]= 7'h0;
assign r_ram[1973]= 7'h0;
assign r_ram[1974]= 7'h49;
assign r_ram[1975]= 7'h0;
assign r_ram[1976]= 7'h0;
assign r_ram[1977]= 7'h0;
assign r_ram[1978]= 7'h0;
assign r_ram[1979]= 7'h0;
assign r_ram[1980]= 7'h0;
assign r_ram[1981]= 7'h0;
assign r_ram[1982]= 7'h0;
assign r_ram[1983]= 7'h0;
assign r_ram[1984]= 7'h4;
assign r_ram[1985]= 7'h0;
assign r_ram[1986]= 7'h8;
assign r_ram[1987]= 7'h0;
assign r_ram[1988]= 7'h0;
assign r_ram[1989]= 7'h0;
assign r_ram[1990]= 7'h0;
assign r_ram[1991]= 7'h2;
assign r_ram[1992]= 7'h0;
assign r_ram[1993]= 7'h0;
assign r_ram[1994]= 7'h0;
assign r_ram[1995]= 7'h0;
assign r_ram[1996]= 7'h0;
assign r_ram[1997]= 7'h0;
assign r_ram[1998]= 7'h0;
assign r_ram[1999]= 7'h0;
assign r_ram[2000]= 7'h0;
assign r_ram[2001]= 7'h0;
assign r_ram[2002]= 7'h11;
assign r_ram[2003]= 7'h0;
assign r_ram[2004]= 7'h0;
assign r_ram[2005]= 7'h0;
assign r_ram[2006]= 7'h0;
assign r_ram[2007]= 7'h0;
assign r_ram[2008]= 7'h0;
assign r_ram[2009]= 7'h0;
assign r_ram[2010]= 7'h0;
assign r_ram[2011]= 7'h0;
assign r_ram[2012]= 7'h0;
assign r_ram[2013]= 7'h0;
assign r_ram[2014]= 7'h0;
assign r_ram[2015]= 7'h0;
assign r_ram[2016]= 7'h0;
assign r_ram[2017]= 7'h0;
assign r_ram[2018]= 7'h0;
assign r_ram[2019]= 7'h0;
assign r_ram[2020]= 7'h2;
assign r_ram[2021]= 7'h0;
assign r_ram[2022]= 7'h0;
assign r_ram[2023]= 7'h0;
assign r_ram[2024]= 7'h0;
assign r_ram[2025]= 7'h0;
assign r_ram[2026]= 7'h0;
assign r_ram[2027]= 7'h0;
assign r_ram[2028]= 7'h0;
assign r_ram[2029]= 7'hc;
assign r_ram[2030]= 7'h0;
assign r_ram[2031]= 7'h0;
assign r_ram[2032]= 7'h0;
assign r_ram[2033]= 7'h0;
assign r_ram[2034]= 7'h0;
assign r_ram[2035]= 7'h0;
assign r_ram[2036]= 7'h21;
assign r_ram[2037]= 7'h0;
assign r_ram[2038]= 7'h0;
assign r_ram[2039]= 7'h0;
assign r_ram[2040]= 7'h0;
assign r_ram[2041]= 7'h0;
assign r_ram[2042]= 7'h0;
assign r_ram[2043]= 7'h0;
assign r_ram[2044]= 7'h0;
assign r_ram[2045]= 7'h0;
assign r_ram[2046]= 7'h0;
assign r_ram[2047]= 7'h0;
assign r_ram[2048]= 7'h0;
assign r_ram[2049]= 7'h0;
assign r_ram[2050]= 7'h2;
assign r_ram[2051]= 7'h0;
assign r_ram[2052]= 7'h0;
assign r_ram[2053]= 7'h0;
assign r_ram[2054]= 7'h0;
assign r_ram[2055]= 7'h0;
assign r_ram[2056]= 7'h0;
assign r_ram[2057]= 7'h0;
assign r_ram[2058]= 7'h0;
assign r_ram[2059]= 7'h0;
assign r_ram[2060]= 7'h0;
assign r_ram[2061]= 7'h0;
assign r_ram[2062]= 7'h0;
assign r_ram[2063]= 7'h0;
assign r_ram[2064]= 7'h8;
assign r_ram[2065]= 7'h4;
assign r_ram[2066]= 7'h0;
assign r_ram[2067]= 7'h0;
assign r_ram[2068]= 7'h41;
assign r_ram[2069]= 7'h0;
assign r_ram[2070]= 7'h0;
assign r_ram[2071]= 7'h0;
assign r_ram[2072]= 7'h0;
assign r_ram[2073]= 7'h0;
assign r_ram[2074]= 7'h0;
assign r_ram[2075]= 7'h0;
assign r_ram[2076]= 7'h4;
assign r_ram[2077]= 7'h0;
assign r_ram[2078]= 7'h0;
assign r_ram[2079]= 7'h8;
assign r_ram[2080]= 7'h0;
assign r_ram[2081]= 7'h2;
assign r_ram[2082]= 7'h0;
assign r_ram[2083]= 7'h0;
assign r_ram[2084]= 7'h0;
assign r_ram[2085]= 7'h0;
assign r_ram[2086]= 7'h0;
assign r_ram[2087]= 7'h0;
assign r_ram[2088]= 7'h0;
assign r_ram[2089]= 7'h0;
assign r_ram[2090]= 7'h0;
assign r_ram[2091]= 7'h0;
assign r_ram[2092]= 7'h0;
assign r_ram[2093]= 7'h11;
assign r_ram[2094]= 7'h0;
assign r_ram[2095]= 7'h0;
assign r_ram[2096]= 7'h0;
assign r_ram[2097]= 7'h0;
assign r_ram[2098]= 7'h0;
assign r_ram[2099]= 7'h0;
assign r_ram[2100]= 7'h0;
assign r_ram[2101]= 7'h0;
assign r_ram[2102]= 7'h0;
assign r_ram[2103]= 7'h0;
assign r_ram[2104]= 7'h0;
assign r_ram[2105]= 7'h0;
assign r_ram[2106]= 7'h0;
assign r_ram[2107]= 7'h0;
assign r_ram[2108]= 7'h0;
assign r_ram[2109]= 7'h0;
assign r_ram[2110]= 7'h2;
assign r_ram[2111]= 7'h0;
assign r_ram[2112]= 7'h0;
assign r_ram[2113]= 7'h0;
assign r_ram[2114]= 7'h0;
assign r_ram[2115]= 7'h0;
assign r_ram[2116]= 7'h8;
assign r_ram[2117]= 7'h0;
assign r_ram[2118]= 7'h4;
assign r_ram[2119]= 7'h0;
assign r_ram[2120]= 7'h0;
assign r_ram[2121]= 7'h0;
assign r_ram[2122]= 7'h0;
assign r_ram[2123]= 7'h0;
assign r_ram[2124]= 7'h0;
assign r_ram[2125]= 7'h21;
assign r_ram[2126]= 7'h0;
assign r_ram[2127]= 7'h0;
assign r_ram[2128]= 7'h0;
assign r_ram[2129]= 7'h0;
assign r_ram[2130]= 7'h0;
assign r_ram[2131]= 7'h0;
assign r_ram[2132]= 7'h0;
assign r_ram[2133]= 7'h0;
assign r_ram[2134]= 7'h0;
assign r_ram[2135]= 7'h0;
assign r_ram[2136]= 7'h0;
assign r_ram[2137]= 7'h0;
assign r_ram[2138]= 7'h0;
assign r_ram[2139]= 7'h0;
assign r_ram[2140]= 7'h2;
assign r_ram[2141]= 7'h0;
assign r_ram[2142]= 7'h0;
assign r_ram[2143]= 7'h0;
assign r_ram[2144]= 7'h0;
assign r_ram[2145]= 7'h0;
assign r_ram[2146]= 7'h0;
assign r_ram[2147]= 7'h0;
assign r_ram[2148]= 7'h0;
assign r_ram[2149]= 7'h4;
assign r_ram[2150]= 7'h0;
assign r_ram[2151]= 7'h0;
assign r_ram[2152]= 7'h8;
assign r_ram[2153]= 7'h0;
assign r_ram[2154]= 7'h0;
assign r_ram[2155]= 7'h0;
assign r_ram[2156]= 7'h41;
assign r_ram[2157]= 7'h0;
assign r_ram[2158]= 7'h0;
assign r_ram[2159]= 7'h0;
assign r_ram[2160]= 7'h0;
assign r_ram[2161]= 7'h0;
assign r_ram[2162]= 7'h0;
assign r_ram[2163]= 7'h0;
assign r_ram[2164]= 7'h0;
assign r_ram[2165]= 7'h0;
assign r_ram[2166]= 7'h8;
assign r_ram[2167]= 7'h4;
assign r_ram[2168]= 7'h0;
assign r_ram[2169]= 7'h0;
assign r_ram[2170]= 7'h0;
assign r_ram[2171]= 7'h2;
assign r_ram[2172]= 7'h0;
assign r_ram[2173]= 7'h0;
assign r_ram[2174]= 7'h0;
assign r_ram[2175]= 7'h0;
assign r_ram[2176]= 7'h0;
assign r_ram[2177]= 7'h0;
assign r_ram[2178]= 7'h0;
assign r_ram[2179]= 7'h0;
assign r_ram[2180]= 7'h0;
assign r_ram[2181]= 7'h0;
assign r_ram[2182]= 7'h0;
assign r_ram[2183]= 7'h11;
assign r_ram[2184]= 7'h0;
assign r_ram[2185]= 7'h0;
assign r_ram[2186]= 7'h0;
assign r_ram[2187]= 7'h0;
assign r_ram[2188]= 7'h0;
assign r_ram[2189]= 7'h0;
assign r_ram[2190]= 7'h0;
assign r_ram[2191]= 7'h0;
assign r_ram[2192]= 7'h0;
assign r_ram[2193]= 7'h0;
assign r_ram[2194]= 7'h0;
assign r_ram[2195]= 7'h0;
assign r_ram[2196]= 7'h0;
assign r_ram[2197]= 7'h0;
assign r_ram[2198]= 7'h0;
assign r_ram[2199]= 7'h0;
assign r_ram[2200]= 7'h2;
assign r_ram[2201]= 7'h0;
assign r_ram[2202]= 7'h0;
assign r_ram[2203]= 7'h0;
assign r_ram[2204]= 7'h0;
assign r_ram[2205]= 7'h0;
assign r_ram[2206]= 7'h4;
assign r_ram[2207]= 7'h8;
assign r_ram[2208]= 7'h0;
assign r_ram[2209]= 7'h0;
assign r_ram[2210]= 7'h0;
assign r_ram[2211]= 7'h0;
assign r_ram[2212]= 7'h0;
assign r_ram[2213]= 7'h0;
assign r_ram[2214]= 7'h0;
assign r_ram[2215]= 7'h0;
assign r_ram[2216]= 7'h21;
assign r_ram[2217]= 7'h0;
assign r_ram[2218]= 7'h0;
assign r_ram[2219]= 7'h0;
assign r_ram[2220]= 7'h0;
assign r_ram[2221]= 7'h0;
assign r_ram[2222]= 7'h0;
assign r_ram[2223]= 7'h0;
assign r_ram[2224]= 7'h0;
assign r_ram[2225]= 7'h0;
assign r_ram[2226]= 7'h0;
assign r_ram[2227]= 7'h0;
assign r_ram[2228]= 7'h0;
assign r_ram[2229]= 7'h0;
assign r_ram[2230]= 7'h0;
assign r_ram[2231]= 7'h2;
assign r_ram[2232]= 7'h0;
assign r_ram[2233]= 7'h0;
assign r_ram[2234]= 7'h0;
assign r_ram[2235]= 7'h0;
assign r_ram[2236]= 7'h0;
assign r_ram[2237]= 7'h0;
assign r_ram[2238]= 7'h0;
assign r_ram[2239]= 7'h0;
assign r_ram[2240]= 7'h0;
assign r_ram[2241]= 7'h0;
assign r_ram[2242]= 7'h4;
assign r_ram[2243]= 7'h0;
assign r_ram[2244]= 7'h0;
assign r_ram[2245]= 7'h8;
assign r_ram[2246]= 7'h41;
assign r_ram[2247]= 7'h0;
assign r_ram[2248]= 7'h0;
assign r_ram[2249]= 7'h0;

endmodule